.model             jjmod                     jj(Rtype=1,  Vg=2.8mV,    Cap=0.064pF,  R0=100ohm,  Rn=17ohm,      Icrit=0.1mA)


.subckt            boost2_4_f4               1            2            3             54          55             56                     57    58    59
*inst name         cell_name                 a            din          dout          q1          q2             q3                     q4    xin   xout
B1                 15                        0            jjmod        area=0.5
B1a                51                        0            jjmod        area=0.5
B1b                19                        0            jjmod        area=0.5
B1c                22                        0            jjmod        area=0.5
B1d                30                        0            jjmod        area=0.5
B2                 34                        0            jjmod        area=0.5
B2a                18                        0            jjmod        area=0.5
B2b                9                         0            jjmod        area=0.5
B2c                20                        0            jjmod        area=0.5
B2d                28                        0            jjmod        area=0.5
Kd1                Ld                        L1           -0.133
Kd1a               Lda                       L1a          -0.133
Kd1b               Ldb                       L1b          -0.133
Kd1c               Ldc                       L1c          -0.133
Kd1d               Ldd                       L1d          -0.133
Kd2                Ld                        L2           -0.133
Kd2a               Lda                       L2a          -0.133
Kd2b               Ldb                       L2b          -0.133
Kd2c               Ldc                       L2c          -0.133
Kd2d               Ldd                       L2d          -0.133
Kdouta             Lda                       Louta        0.0
Kdoutb             Ldb                       Loutb        0.0
Kdoutc             Ldc                       Loutc        0.0
Kdoutd             Ldd                       Loutd        0.0
Kdqa               Lda                       Lqa          0.0
Kdqb               Ldb                       Lqb          0.0
Kdqc               Ldc                       Lqc          0.0
Kdqd               Ldd                       Lqd          0.0
Kouta              Lqa                       Louta        -0.495
Koutb              Lqb                       Loutb        -0.495
Koutd              Lqd                       Loutd        -0.495
Kqoutc             Lqc                       Loutc        -0.495
Kx1                Lx                        L1           -0.186
Kx1a               Lxa                       L1a          -0.186
Kx1b               Lxb                       L1b          -0.186
Kx1c               Lxc                       L1c          -0.186
Kx1d               Lxd                       L1d          -0.186
Kx2                Lx                        L2           -0.186
Kx2a               Lxa                       L2a          -0.186
Kx2b               Lxb                       L2b          -0.186
Kx2c               Lxc                       L2c          -0.186
Kx2d               Lxd                       L2d          -0.186
Kxd                Lx                        Ld           0.19
Kxda               Lxa                       Lda          0.19
Kxdb               Lxb                       Ldb          0.19
Kxdc               Lxc                       Ldc          0.19
Kxdd               Lxd                       Ldd          0.19
Kxouta             Lxa                       Louta        0.0
Kxoutb             Lxb                       Loutb        0.0
Kxoutc             Lxc                       Loutc        0.0
Kxoutd             Lxd                       Loutd        0.0
Kxqa               Lxa                       Lqa          0.0
Kxqb               Lxb                       Lqb          0.0
Kxqc               Lxc                       Lqc          0.0
Kxqd               Lxd                       Lqd          0.0
L1                 45                        15           1.59pH
L1a                50                        51           1.59pH
L1b                49                        19           1.59pH
L1c                40                        22           1.59pH
L1d                48                        30           1.59pH
L2                 34                        45           1.59pH
L2a                18                        50           1.59pH
L2b                9                         49           1.59pH
L2c                20                        40           1.59pH
L2d                28                        48           1.59pH
Ld                 2                         6            7.45pH
Lda                6                         5            7.45pH
Ldb                5                         41           7.45pH
Ldc                41                        46           7.45pH
Ldd                46                        3            7.45pH
Lin                1                         45           1.23pH
Lina               4                         50           3.4pH
Linb               4                         49           3.0pH
Linc               4                         40           3.0pH
Lind               4                         48           3.4pH
Louta              25                        54           31.2pH
Loutb              17                        55           31.2pH
Loutc              38                        56           31.2pH
Loutd              47                        57           31.2pH
Lq                 45                        4            9.96pH
Lqa                50                        53           7.92pH
Lqb                49                        24           7.92pH
Lqc                40                        26           7.92pH
Lqd                48                        32           7.92pH
Lx                 58                        7            7.4pH
Lxa                7                         8            7.4pH
Lxb                8                         16           7.4pH
Lxc                16                        43           7.4pH
Lxd                43                        59           7.4pH
R1a                25                        0            1e-12ohm
R1b                17                        0            1e-12ohm
R4                 53                        0            1e-12ohm
R5                 24                        0            1e-12ohm
R6                 38                        0            1e-12ohm
R7                 26                        0            1e-12ohm
R8                 47                        0            1e-12ohm
R9                 32                        0            1e-12ohm
.ends


.subckt            branch3                   1            2            3             4
*inst name         cell_name                 a            b            c             d
Lip                7                         4            0.312pH
Lp1                1                         6            11.8pH
Lp2                2                         7            10.2pH
Lp3                3                         5            11.8pH
R0                 6                         7            1e-12ohm
R1                 5                         7            1e-12ohm
.ends


.subckt            const0                    1            2            11            12          13
*inst name         cell_name                 din          dout         q             xin         xout
B1                 8                         0            jjmod        area=0.5
B2                 4                         0            jjmod        area=0.5
Kd1                Ld                        L1           -0.128
Kd2                Ld                        L2           -0.135
Kdout              Ld                        Lout         -0.000253
Kdq                Ld                        Lq           -0.00468
Kout               Lq                        Lout         -0.495
Kx1                Lx                        L1           -0.185
Kx2                Lx                        L2           -0.189
Kxd                Lx                        Ld           0.193
Kxout              Lx                        Lout         -7.94e-05
Kxq                Lx                        Lq           -0.00421
L1                 7                         8            1.56pH
L2                 4                         7            1.66pH
Ld                 1                         2            7.49pH
Lout               5                         11           31.2pH
Lq                 7                         0            7.82pH
Lx                 12                        13           7.47pH
R1                 5                         0            1e-12ohm
.ends


.subckt            bfr                       1            2            3             12          13             14
*inst name         cell_name                 a            din          dout          q           xin            xout
B1                 9                         0            jjmod        area=0.5
B2                 5                         0            jjmod        area=0.5
Kd1                Ld                        L1           -0.133
Kd2                Ld                        L2           -0.133
Kdout              Ld                        Lout         0.0
Kdq                Ld                        Lq           0.0
Kout               Lq                        Lout         -0.495
Kx1                Lx                        L1           -0.186
Kx2                Lx                        L2           -0.186
Kxd                Lx                        Ld           0.19
Kxout              Lx                        Lout         0.0
Kxq                Lx                        Lq           0.0
L1                 8                         9            1.59pH
L2                 5                         8            1.59pH
Ld                 2                         3            7.45pH
Lin                1                         8            1.23pH
Lout               6                         12           31.2pH
Lq                 8                         0            7.92pH
Lx                 13                        14           7.4pH
R1                 6                         0            1e-12ohm
.ends


.subckt            and_bb                    1            2            3             4           12             13                     14
*inst name         cell_name                 a            b            din           dout        q              xin                    xout
XI0                bfr                       1            3            8             9           13             5
XI2                bfr                       2            11           4             10          7              14
XI3                branch3                   9            6            10            12
XI1                const0                    8            11           6             5           7
.ends


.subckt            inv                       1            2            3             12          13             14
*inst name         cell_name                 a            din          dout          q           xin            xout
B1                 9                         0            jjmod        area=0.6
B2                 5                         0            jjmod        area=0.6
Kd1                Ld                        L1           -0.133
Kd2                Ld                        L2           -0.133
Kdout              Ld                        Lout         0.0
Kdq                Ld                        Lq           0.0
Kout               Lq                        Lout         0.432
Kx1                Lx                        L1           -0.186
Kx2                Lx                        L2           -0.186
Kxd                Lx                        Ld           0.19
Kxout              Lx                        Lout         0.0
Kxq                Lx                        Lq           0.0
L1                 8                         9            1.59pH
L2                 5                         8            1.59pH
Ld                 2                         3            7.44pH
Lin                1                         8            1.24pH
Lout               6                         12           31.0pH
Lq                 8                         0            6.49pH
Lx                 13                        14           7.39pH
R1                 6                         0            1e-12ohm
.ends


.subckt            maj_bbi                   1            2            3             4           5              13                     14    15
*inst name         cell_name                 a            b            c             din         dout           q                      xin   xout
XI0                bfr                       1            4            9             11          14             6
XI1                bfr                       2            9            12            7           6              8
XI3                branch3                   11           7            10            13
XI2                inv                       3            12           5             10          8              15
.ends


.subckt            boost2_3_f3               1            2            3             41          42             43                     44    45
*inst name         cell_name                 a            din          dout          q1          q2             q3                     xin   xout
B1                 11                        0            jjmod        area=0.5
B1a                36                        0            jjmod        area=0.5
B1b                14                        0            jjmod        area=0.5
B1c                17                        0            jjmod        area=0.5
B2                 24                        0            jjmod        area=0.5
B2a                13                        0            jjmod        area=0.5
B2b                5                         0            jjmod        area=0.5
B2c                15                        0            jjmod        area=0.5
Kd1                Ld                        L1           -0.0644
Kd1a               Ld                        L1a          -0.0639
Kd1b               Ld                        L1b          -0.0662
Kd1c               Ld                        L1c          -0.066
Kd2                Ld                        L2           -0.0646
Kd2a               Ld                        L2a          -0.0653
Kd2b               Ld                        L2b          -0.0666
Kd2c               Ld                        L2c          -0.0642
Kdouta             Ld                        Louta        0.0007254
Kdoutb             Ld                        Loutb        0.0004117
Kdoutc             Ld                        Loutc        -0.001253
Kdq                Ld                        Lq           0.0
Kdqa               Ld                        Lqa          -0.0006276
Kdqb               Ld                        Lqb          -0.0005469
Kdqc               Ld                        Lqc          0.001507
Kdql               Ld                        Lql          0.0
Kdqr               Ld                        Lqr          0.0
Kouta              Lqa                       Louta        -0.493
Koutb              Lqb                       Loutb        -0.493
Koutc              Lqc                       Loutc        -0.493
Kx1                Lx                        L1           -0.0881
Kx1a               Lx                        L1a          -0.0893
Kx1b               Lx                        L1b          -0.0909
Kx1c               Lx                        L1c          -0.0907
Kx2                Lx                        L2           -0.0885
Kx2a               Lx                        L2a          -0.0903
Kx2b               Lx                        L2b          -0.0908
Kx2c               Lx                        L2c          -0.0894
Kxd                Lx                        Ld           0.177
Kxouta             Lx                        Louta        0.0003079
Kxoutb             Lx                        Loutb        -9.704e-05
Kxoutc             Lx                        Loutc        -0.0003689
Kxq                Lx                        Lq           0.0
Kxqa               Lx                        Lqa          -0.0003187
Kxqb               Lx                        Lqb          -0.0003226
Kxqc               Lx                        Lqc          0.0008805
Kxql               Lx                        Lql          0.0
Kxqr               Lx                        Lqr          0.0
L1                 31                        11           1.58pH
L1a                34                        36           1.49pH
L1b                32                        14           1.49pH
L1c                29                        17           1.49pH
L2                 24                        31           1.58pH
L2a                13                        34           1.49pH
L2b                5                         32           1.49pH
L2c                15                        29           1.49pH
Ld                 2                         3            36.97pH
Lin                1                         31           2.03pH
Lina               33                        34           1.23pH
Linb               4                         32           1.37pH
Linc               37                        29           1.36pH
Louta              20                        41           31.1pH
Loutb              12                        42           31.1pH
Loutc              27                        43           31.1pH
Lq                 31                        35           7.76pH
Lqa                34                        39           7.9pH
Lqb                32                        19           7.89pH
Lqc                29                        21           7.91pH
Lql                35                        33           5.27pH
Lqr                40                        35           5.06pH
Lqrb               40                        4            0.19pH
Lqrc               40                        37           1.36pH
Lx                 44                        45           36.64pH
R1a                20                        0            1e-12ohm
R1b                12                        0            1e-12ohm
R4                 39                        0            1e-12ohm
R5                 19                        0            1e-12ohm
R6                 27                        0            1e-12ohm
R7                 21                        0            1e-12ohm
.ends


.subckt            maj_bib                   1            2            3             4           5              13                     14    15
*inst name         cell_name                 a            b            c             din         dout           q                      xin   xout
XI0                bfr                       1            4            9             11          14             6
XI2                bfr                       3            7            5             10          8              15
XI3                branch3                   11           12           10            13
XI1                inv                       2            9            7             12          6              8
.ends


.subckt            maj_ibb                   1            2            3             4           5              13                     14    15
*inst name         cell_name                 a            b            c             din         dout           q                      xin   xout
XI1                bfr                       2            8            10            12          6              7
XI2                bfr                       3            10           5             9           7              15
XI3                branch3                   11           12           9             13
XI0                inv                       1            4            8             11          14             6
.ends


.subckt            maj_bbb                   1            2            3             4           5              13                     14    15
*inst name         cell_name                 a            b            c             din         dout           q                      xin   xout
XI0                bfr                       1            4            8             11          14             6
XI1                bfr                       2            8            10            12          6              7
XI2                bfr                       3            10           5             9           7              15
XI3                branch3                   11           12           9             13
.ends


.subckt            sink                      1            2            3             10          11
*inst name         cell_name                 a            din          dout          xin         xout
B1                 8                         0            jjmod        area=0.5
B2                 5                         0            jjmod        area=0.5
Kd1                Ld                        L1           -0.133
Kd2                Ld                        L2           -0.133
Kdq                Ld                        Lq           0.0
Kx1                Lx                        L1           -0.186
Kx2                Lx                        L2           -0.186
Kxd                Lx                        Ld           0.19
Kxq                Lx                        Lq           0.0
L1                 7                         8            1.59pH
L2                 5                         7            1.59pH
Ld                 2                         3            7.45pH
Lin                1                         7            1.23pH
Lq                 7                         0            7.92pH
Lx                 10                        11           7.4pH
.ends


.subckt            and_bi                    1            2            3             4           12             13                     14
*inst name         cell_name                 a            b            din           dout        q              xin                    xout
XI0                bfr                       1            3            8             9           13             5
XI3                branch3                   9            7            10            12
XI1                const0                    8            11           7             5           6
XI2                inv                       2            11           4             10          6              14
.ends


.subckt            and_ib                    1            2            3             4           12             13                     14
*inst name         cell_name                 a            b            din           dout        q              xin                    xout
XI2                bfr                       2            11           4             10          6              14
XI3                branch3                   9            8            10            12
XI1                const0                    7            11           8             5           6
XI0                inv                       1            3            7             9           13             5
.ends


.subckt            const1                    1            2            7             8           9
*inst name         cell_name                 din          dout         q             xin         xout
L1                 8                         4            0.01pH
L2                 6                         9            0.01pH
L3                 1                         3            0.01pH
L4                 5                         2            0.01pH
XI0                const0                    5            3            7             6           4
.ends


.subckt            or_bb                     1            2            3             4           12             13                     14
*inst name         cell_name                 a            b            din           dout        q              xin                    xout
XI0                bfr                       1            3            8             9           13             5
XI2                bfr                       2            11           4             10          6              14
XI3                branch3                   9            7            10            12
XI1                const1                    8            11           7             5           6
.ends


*this is top cell  4bit_RCA_ene_opt_booster
R10                259                       373          1000.0ohm
R3                 265                       357          1000.0ohm
R4                 248                       279          1000.0ohm
R5                 245                       167          1000.0ohm
R6                 249                       171          1000.0ohm
R7                 255                       363          1000.0ohm
R8                 186                       382          1000.0ohm
R9                 182                       347          1000.0ohm
Rac1               253                       413          100000.0ohm
Rac2               240                       416          100000.0ohm
Rdc1               269                       80           100000.0ohm
V10                259                       0            PWL          (0ps          0mv  20ps           {{input[0]}})
V2                 265                       0            PWL          (0ps          0mv 20ps           {{input[1]}})
V4                 248                       0            PWL          (0ps          0mv 20ps           {{input[2]}})
V5                 245                       0            PWL          (0ps          0mv 20ps           {{input[3]}})
V6                 249                       0            PWL          (0ps          0mv 20ps           {{input[4]}})
V7                 255                       0            PWL          (0ps          0mv 20ps           {{input[5]}})
V8                 186                       0            PWL          (0ps          0mv 20ps           {{input[6]}})
V9                 182                       0            PWL          (0ps          0mv 20ps           {{input[7]}})
VDC                269                       0            PWL          (0ps          0mV         20ps           113000mV)
VAC1               253                       0            SIN          (0            81000mV     {{freq}}MEGHz  {{40+period|int/4}}ps  0)
VAC2               240                       0            SIN          (0            81000mV     {{freq}}MEGHz  40ps                   0)
XI333              and_bb                    212          183          73            197         175            124                    76
XI336              and_bi                    161          189          158           73          184            400                    124
XI338              and_ib                    195          194          173           158         215            122                    400
XI100              bfr                       309          341          154           372         209            153
XI101              bfr                       16           288          341           67          285            209
XI102              bfr                       354          322          288           360         412            285
XI103              bfr                       316          369          203           18          219            202
XI104              bfr                       364          214          369           33          281            219
XI105              bfr                       304          216          214           323         346            281
XI106              bfr                       27           198          216           309         328            346
XI107              bfr                       385          386          198           16          333            328
XI108              bfr                       365          322          386           354         416            333
XI109              bfr                       297          326          371           7           338            152
XI110              bfr                       30           286          326           13          344            338
XI111              bfr                       31           351          286           94          208            344
XI112              bfr                       372          205          351           2           207            208
XI113              bfr                       67           355          205           19          290            207
XI114              bfr                       360          243          355           28          415            290
XI117              bfr                       406          314          292           105         83             164
XI118              bfr                       105          230          181           224         69             180
XI119              bfr                       282          292          238           236         164            317
XI120              bfr                       150          264          234           282         329            233
XI121              bfr                       236          181          387           287         180            334
XI122              bfr                       409          310          96            150         370            227
XI123              bfr                       390          238          169           327         317            185
XI124              bfr                       327          387          177           349         334            411
XI125              bfr                       20           96           228           4           227            185
XI126              bfr                       410          232          398           12          391            122
XI127              bfr                       4            234          169           390         233            235
XI128              bfr                       12           84           228           20          401            235
XI129              bfr                       2            193          178           41          191            1
XI130              bfr                       94           178          218           46          1              3
XI131              bfr                       7            176          95            26          5              6
XI132              bfr                       13           218          176           34          3              5
XI133              bfr                       72           179          226           82          239            29
XI134              bfr                       19           221          193           72          166            191
XI135              bfr                       46           22           278           56          211            62
XI136              bfr                       56           37           78            68          23             24
XI137              bfr                       28           243          221           70          412            166
XI138              bfr                       34           278          60            407         62             275
XI139              bfr                       26           60           197           408         275            76
XI140              bfr                       68           274          273           405         272            81
XI141              bfr                       61           256          274           404         39             272
XI142              bfr                       106          74           268           402         54             168
XI143              bfr                       109          268          92            403         168            103
XI144              bfr                       98           47           48            106         49             199
XI145              bfr                       102          48           376           109         199            204
XI146              bfr                       86           47           174           98          54             246
XI147              bfr                       77           36           44            86          49             45
XI148              bfr                       82           44           146           91          45             159
XI149              bfr                       91           174          256           102         246            39
XI150              bfr                       50           146          37            61          159            23
XI151              bfr                       70           36           179           77          415            239
XI152              bfr                       41           226          22            50          29             211
XI332              bfr                       367          138          399           149         0              113
XI59               bfr                       349          90           177           59          88             187
XI60               bfr                       336          117          115           295         110            187
XI61               bfr                       59           119          115           336         112            411
XI63               bfr                       287          108          90            63          125            88
XI64               bfr                       381          100          117           340         99             110
XI65               bfr                       63           308          119           381         130            112
XI67               bfr                       224          296          108           66          101            125
XI68               bfr                       65           104          100           64          141            99
XI69               bfr                       66           378          308           65          128            130
XI71               bfr                       188          192          139           53          395            85
XI72               bfr                       52           111          142           367         107            134
XI73               bfr                       53           111          135           52          414            143
XI75               bfr                       133          135          296           313         143            101
XI76               bfr                       55           399          104           51          113            141
XI77               bfr                       313          142          378           55          134            128
XI83               bfr                       357          299          147           339         289            388
XI84               bfr                       279          301          299           321         397            289
XI85               bfr                       330          379          300           302         311            388
XI86               bfr                       58           244          379           57          120            311
XI87               bfr                       339          280          147           330         306            163
XI88               bfr                       321          203          280           58          202            306
XI89               bfr                       302          267          300           210         362            163
XI90               bfr                       57           371          267           190         152            362
XI91               bfr                       167          201          301           316         342            397
XI92               bfr                       171          361          201           364         229            342
XI93               bfr                       363          380          361           304         172            229
XI94               bfr                       382          318          380           27          271            172
XI95               bfr                       347          359          318           385         276            271
XI96               bfr                       373          80           359           365         413            276
XI97               bfr                       18           396          244           297         384            120
XI98               bfr                       33           148          396           30          374            384
XI99               bfr                       323          154          148           31          153            374
XI340              boost2_3_f3               190          95           127           183         189            194                    6     126
XI341              boost2_3_f3               210          127          173           212         161            195                    126   157
XI312              boost2_4_f4               407          78           320           293         220            206                    196   24    38
XI313              boost2_4_f4               408          320          375           217         213            343                    393   38    394
XI314              boost2_4_f4               175          375          160           200         315            241                    247   394   97
XI316              boost2_4_f4               404          376          25            170         151            155                    145   204   10
XI321              boost2_4_f4               405          25           277           165         156            123                    118   10    21
XI322              boost2_4_f4               324          277          75            136         140            116                    307   21    93
XI323              boost2_4_f4               402          74           35            353         358            356                    392   395   17
XI326              boost2_4_f4               403          35           303           383         348            283                    319   17    11
XI329              boost2_4_f4               298          303          89            332         368            260                    305   11    79
XI307              maj_bbb                   293          217          200           273         350            324                    81    294
XI310              maj_bbb                   325          237          366           75          84             409                    93    401
XI315              maj_bbb                   170          165          136           92          270            298                    103   32
XI318              maj_bbb                   162          291          129           89          264            406                    79    329
XI324              maj_bbb                   353          383          332           192         43             188                    414   15
XI330              maj_bbb                   335          389          284           139         230            133                    85    69
XI311              maj_bbi                   196          393          247           8           232            366                    9     391
XI317              maj_bbi                   145          118          307           345         310            129                    257   370
XI328              maj_bbi                   392          319          305           312         314            284                    337   83
XI309              maj_bib                   206          343          241           377         8              237                    352   9
XI319              maj_bib                   155          123          116           42          345            291                    40    257
XI327              maj_bib                   356          283          260           14          312            389                    331   337
XI308              maj_ibb                   220          213          315           350         377            325                    294   352
XI320              maj_ibb                   151          156          140           270         42             162                    32    40
XI325              maj_ibb                   358          348          368           43          14             335                    15    331
XI339              or_bb                     184          215          160           398         410            97                     157
XSUM0              sink                      295          251          0             114         0
XSUM1              sink                      340          131          251           132         114
XSUM2              sink                      64           254          131           144         132
XSUM3              sink                      51           121          254           137         144
XSUM4              sink                      149          138          121           107         137
*end of top cell   4bit_RCA_ene_opt_booster


.tran              {{t_step}}ps              {{end}}ps    {{begin}}ps  {{t_step}}ps
.FiLE              {{out_file_name}}
.print             i(Rac1)
*vac1_tot
.print             nodev                     413          0

.print             i(Rac2)
*vac2_tot
.print             nodev                     416          0

*vac1_DUT
.print             nodev                     412          411
*vac2_DUT
.print             nodev                     415          414
