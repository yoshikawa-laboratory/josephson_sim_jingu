.model             jjmod                           jj(Rtype=1,  Vg=2.8mV,    Cap=0.064pF,  R0=100ohm,  Rn=17ohm,      Icrit=0.1mA)


.subckt            branch3                         1            2            3             4
*inst name         cell_name                       a            b            c             d
Lip                7                               4            0.312pH
Lp1                1                               6            11.8pH
Lp2                2                               7            10.2pH
Lp3                3                               5            11.8pH
R0                 6                               7            1e-12ohm
R1                 5                               7            1e-12ohm
.ends


.subckt            const0                          1            2            11            12          13
*inst name         cell_name                       din          dout         q             xin         xout
B1                 8                               0            jjmod        area=0.5
B2                 4                               0            jjmod        area=0.5
Kd1                Ld                              L1           -0.128
Kd2                Ld                              L2           -0.135
Kdout              Ld                              Lout         -0.000253
Kdq                Ld                              Lq           -0.00468
Kout               Lq                              Lout         -0.495
Kx1                Lx                              L1           -0.185
Kx2                Lx                              L2           -0.189
Kxd                Lx                              Ld           0.193
Kxout              Lx                              Lout         -7.94e-05
Kxq                Lx                              Lq           -0.00421
L1                 7                               8            1.56pH
L2                 4                               7            1.66pH
Ld                 1                               2            7.49pH
Lout               5                               11           31.2pH
Lq                 7                               0            7.82pH
Lx                 12                              13           7.47pH
R1                 5                               0            1e-12ohm
.ends


.subckt            bfr                             1            2            3             12          13             14
*inst name         cell_name                       a            din          dout          q           xin            xout
B1                 9                               0            jjmod        area=0.5
B2                 5                               0            jjmod        area=0.5
Kd1                Ld                              L1           -0.133
Kd2                Ld                              L2           -0.133
Kdout              Ld                              Lout         0.0
Kdq                Ld                              Lq           0.0
Kout               Lq                              Lout         -0.495
Kx1                Lx                              L1           -0.186
Kx2                Lx                              L2           -0.186
Kxd                Lx                              Ld           0.19
Kxout              Lx                              Lout         0.0
Kxq                Lx                              Lq           0.0
L1                 8                               9            1.59pH
L2                 5                               8            1.59pH
Ld                 2                               3            7.45pH
Lin                1                               8            1.23pH
Lout               6                               12           31.2pH
Lq                 8                               0            7.92pH
Lx                 13                              14           7.4pH
R1                 6                               0            1e-12ohm
.ends


.subckt            and_bb                          1            2            3             4           12             13                     14
*inst name         cell_name                       a            b            din           dout        q              xin                    xout
XI0                bfr                             1            3            8             9           13             5
XI2                bfr                             2            11           4             10          7              14
XI3                branch3                         9            6            10            12
XI1                const0                          8            11           6             5           7
.ends


.subckt            const1                          1            2            7             8           9
*inst name         cell_name                       din          dout         q             xin         xout
L1                 8                               4            0.01pH
L2                 6                               9            0.01pH
L3                 1                               3            0.01pH
L4                 5                               2            0.01pH
XI0                const0                          5            3            7             6           4
.ends


.subckt            or_bb                           1            2            3             4           12             13                     14
*inst name         cell_name                       a            b            din           dout        q              xin                    xout
XI0                bfr                             1            3            8             9           13             5
XI2                bfr                             2            11           4             10          6              14
XI3                branch3                         9            7            10            12
XI1                const1                          8            11           7             5           6
.ends


.subckt            bias_pair_10um                  1            2            3             4
*inst name         cell_name                       a            b            c             d
*C0                 2                               0            0.00145pF
*C6                 4                               0            0.00144pF
L0                 1                               2            3.46pH
L1                 3                               4            3.73pH
.ends


.subckt            branch2                         1            2            3
*inst name         cell_name                       a            b            c
Lip                6                               3            0.282pH
Lp1                1                               5            11.0pH
Lp2                2                               4            11.0pH
R0                 5                               6            1e-12ohm
R1                 4                               6            1e-12ohm
.ends


.subckt            spl2                            1            2            3             9           10             11                     12
*inst name         cell_name                       a            din          dout          x           xin            xout                   y
XI0                bfr                             1            4            6             7           8              5
XI14               bias_pair_10um                  10           8            2             4
XI15               bias_pair_10um                  5            11           6             3
XI1                branch2                         9            12           7
.ends


.subckt            maj_bbb                         1            2            3             4           5              13                     14         15
*inst name         cell_name                       a            b            c             din         dout           q                      xin        xout
XI0                bfr                             1            4            8             11          14             6
XI1                bfr                             2            8            10            12          6              7
XI2                bfr                             3            10           5             9           7              15
XI3                branch3                         11           12           9             13
.ends


.subckt            boost2_3_f3                     1            2            3             41          42             43                     44         45
*inst name         cell_name                       a            din          dout          q1          q2             q3                     xin        xout
B1                 11                              0            jjmod        area=0.5
B1a                36                              0            jjmod        area=0.5
B1b                14                              0            jjmod        area=0.5
B1c                17                              0            jjmod        area=0.5
B2                 24                              0            jjmod        area=0.5
B2a                13                              0            jjmod        area=0.5
B2b                5                               0            jjmod        area=0.5
B2c                15                              0            jjmod        area=0.5
Kd1                Ld                              L1           -0.0644
Kd1a               Ld                              L1a          -0.0639
Kd1b               Ld                              L1b          -0.0662
Kd1c               Ld                              L1c          -0.066
Kd2                Ld                              L2           -0.0646
Kd2a               Ld                              L2a          -0.0653
Kd2b               Ld                              L2b          -0.0666
Kd2c               Ld                              L2c          -0.0642
Kdouta             Ld                              Louta        0.0007254
Kdoutb             Ld                              Loutb        0.0004117
Kdoutc             Ld                              Loutc        -0.001253
Kdq                Ld                              Lq           0.0
Kdqa               Ld                              Lqa          -0.0006276
Kdqb               Ld                              Lqb          -0.0005469
Kdqc               Ld                              Lqc          0.001507
Kdql               Ld                              Lql          0.0
Kdqr               Ld                              Lqr          0.0
Kouta              Lqa                             Louta        -0.493
Koutb              Lqb                             Loutb        -0.493
Koutc              Lqc                             Loutc        -0.493
Kx1                Lx                              L1           -0.0881
Kx1a               Lx                              L1a          -0.0893
Kx1b               Lx                              L1b          -0.0909
Kx1c               Lx                              L1c          -0.0907
Kx2                Lx                              L2           -0.0885
Kx2a               Lx                              L2a          -0.0903
Kx2b               Lx                              L2b          -0.0908
Kx2c               Lx                              L2c          -0.0894
Kxd                Lx                              Ld           0.177
Kxouta             Lx                              Louta        0.0003079
Kxoutb             Lx                              Loutb        -9.704e-05
Kxoutc             Lx                              Loutc        -0.0003689
Kxq                Lx                              Lq           0.0
Kxqa               Lx                              Lqa          -0.0003187
Kxqb               Lx                              Lqb          -0.0003226
Kxqc               Lx                              Lqc          0.0008805
Kxql               Lx                              Lql          0.0
Kxqr               Lx                              Lqr          0.0
L1                 31                              11           1.58pH
L1a                34                              36           1.49pH
L1b                32                              14           1.49pH
L1c                29                              17           1.49pH
L2                 24                              31           1.58pH
L2a                13                              34           1.49pH
L2b                5                               32           1.49pH
L2c                15                              29           1.49pH
Ld                 2                               3            36.97pH
Lin                1                               31           2.03pH
Lina               33                              34           1.23pH
Linb               4                               32           1.37pH
Linc               37                              29           1.36pH
Louta              20                              41           31.1pH
Loutb              12                              42           31.1pH
Loutc              27                              43           31.1pH
Lq                 31                              35           7.76pH
Lqa                34                              39           7.9pH
Lqb                32                              19           7.89pH
Lqc                29                              21           7.91pH
Lql                35                              33           5.27pH
Lqr                40                              35           5.06pH
Lqrb               40                              4            0.19pH
Lqrc               40                              37           1.36pH
Lx                 44                              45           36.64pH
R1a                20                              0            1e-12ohm
R1b                12                              0            1e-12ohm
R4                 39                              0            1e-12ohm
R5                 19                              0            1e-12ohm
R6                 27                              0            1e-12ohm
R7                 21                              0            1e-12ohm
.ends


.subckt            inv                             1            2            3             12          13             14
*inst name         cell_name                       a            din          dout          q           xin            xout
B1                 9                               0            jjmod        area=0.6
B2                 5                               0            jjmod        area=0.6
Kd1                Ld                              L1           -0.133
Kd2                Ld                              L2           -0.133
Kdout              Ld                              Lout         0.0
Kdq                Ld                              Lq           0.0
Kout               Lq                              Lout         0.432
Kx1                Lx                              L1           -0.186
Kx2                Lx                              L2           -0.186
Kxd                Lx                              Ld           0.19
Kxout              Lx                              Lout         0.0
Kxq                Lx                              Lq           0.0
L1                 8                               9            1.59pH
L2                 5                               8            1.59pH
Ld                 2                               3            7.44pH
Lin                1                               8            1.24pH
Lout               6                               12           31.0pH
Lq                 8                               0            6.49pH
Lx                 13                              14           7.39pH
R1                 6                               0            1e-12ohm
.ends


.subckt            maj_bbi                         1            2            3             4           5              13                     14         15
*inst name         cell_name                       a            b            c             din         dout           q                      xin        xout
XI0                bfr                             1            4            9             11          14             6
XI1                bfr                             2            9            12            7           6              8
XI3                branch3                         11           7            10            13
XI2                inv                             3            12           5             10          8              15
.ends


.subckt            maj_ibb                         1            2            3             4           5              13                     14         15
*inst name         cell_name                       a            b            c             din         dout           q                      xin        xout
XI1                bfr                             2            8            10            12          6              7
XI2                bfr                             3            10           5             9           7              15
XI3                branch3                         11           12           9             13
XI0                inv                             1            4            8             11          14             6
.ends


.subckt            maj3_KSA_sum_ene_opt_boost      1            2            3             4           5              6                      7          8     9         10        11         12         13         14         15         34
*inst name         cell_name                       a            ac_in<0>     ac_in<1>      ac_in<2>    ac_out<0>      ac_out<1>              ac_out<2>  b     c         dc_in<0>  dc_in<1>   dc_in<2>   dc_out<0>  dc_out<1>  dc_out<2>  sum
XI3                bfr                             27           30           14            18          29             6
XI18               boost2_3_f3                     9            15           21            27          32             31                     7          20
XI0                maj_bbb                         24           17           31            11          28             33                     3          26
XI1                maj_bbi                         25           23           32            28          30             16                     26         29
XI2                maj_ibb                         33           16           18            10          13             34                     2          5
XI16               spl2                            8            22           21            17          19             20                     23
XI6                spl2                            1            12           22            24          4              19                     25
.ends


.subckt            maj3_KSA_GP_ene_opt             1            2            3             4           5              6                      7          8     9         10        11         12
*inst name         cell_name                       G            P            a             ac_in<0>    ac_in<1>       ac_out<0>              ac_out<1>  b     dc_in<0>  dc_in<1>  dc_out<0>  dc_out<1>
XI9                and_bb                          13           14           19            9           1              20                     4
XI10               or_bb                           18           16           11            19          2              6                      20
XI11               spl2                            3            10           17            14          5              15                     16
XI12               spl2                            8            17           12            13          15             7                      18
.ends


.subckt            sink                            1            2            3             10          11
*inst name         cell_name                       a            din          dout          xin         xout
B1                 8                               0            jjmod        area=0.5
B2                 5                               0            jjmod        area=0.5
Kd1                Ld                              L1           -0.133
Kd2                Ld                              L2           -0.133
Kdq                Ld                              Lq           0.0
Kx1                Lx                              L1           -0.186
Kx2                Lx                              L2           -0.186
Kxd                Lx                              Ld           0.19
Kxq                Lx                              Lq           0.0
L1                 7                               8            1.59pH
L2                 5                               7            1.59pH
Ld                 2                               3            7.45pH
Lin                1                               7            1.23pH
Lq                 7                               0            7.92pH
Lx                 10                              11           7.4pH
.ends


*this is top cell  maj3_4_bit_KSA_ene_opt_booster
R0                 366                             343          1000.0ohm
R1                 363                             373          1000.0ohm
R2                 377                             521          1000.0ohm
R3                 372                             388          1000.0ohm
R4                 369                             181          1000.0ohm
R5                 375                             402          1000.0ohm
R6                 360                             520          1000.0ohm
R7                 359                             357          1000.0ohm
R9                 222                             16           100000.0ohm
Rac1               456                             528          100000.0ohm
Rac2               180                             531          100000.0ohm
V12                366                             0            PWL          (0ps          0mv         20ps           {{input[0]}})
V13                377                             0            PWL          (0ps          0mv         20ps           {{input[1]}})
V14                369                             0            PWL          (0ps          0mv         20ps           {{input[2]}})
V15                360                             0            PWL          (0ps          0mv         20ps           {{input[3]}})
V16                363                             0            PWL          (0ps          0mv         20ps           {{input[4]}})
V17                372                             0            PWL          (0ps          0mv         20ps           {{input[5]}})
V18                375                             0            PWL          (0ps          0mv         20ps           {{input[6]}})
V19                359                             0            PWL          (0ps          0mv         20ps           {{input[7]}})
VDC                222                             0            PWL          (0ps          0mV         20ps           113000mV)
VAC1               456                             0            SIN          (0            81000mV     {{freq}}MEGHz  {{40+period|int/4}}ps  0)
VAC2               180                             0            SIN          (0            81000mV     {{freq}}MEGHz  40ps                   0)
XI1089             and_bb                          187          420          17            524         512            511                    523
XI1092             and_bb                          193          489          497           477         481            510                    470
XI440              and_bb                          271          278          251           289         291            253                    288
XI441              and_bb                          228          286          283           294         296            284                    293
XI1014             bfr                             213          115          111           212         460            112
XI102              bfr                             370          391          315           263         389            314
XI1027             bfr                             236          147          49            218         145            303
XI105              bfr                             252          397          414           384         396            413
XI106              bfr                             507          418          19            301         416            209
XI1090             bfr                             522          519          524           387         518            523
XI1093             bfr                             464          450          477           390         444            470
XI1100             bfr                             513          432          429           514         133            431
XI1101             bfr                             192          129          424           189         371            423
XI1102             bfr                             422          424          428           437         423            425
XI1103             bfr                             198          300          452           196         18             123
XI1113             bfr                             208          452          116           210         123            459
XI1114             bfr                             212          116          113           195         459            114
XI1115             bfr                             217          113          119           149         114            118
XI1116             bfr                             203          206          458           207         205            117
XI1117             bfr                             218          458          100           219         117            101
XI112              bfr                             185          299          172           12          526            161
XI113              bfr                             12           65           66            11          529            67
XI114              bfr                             11           65           64            13          0              175
XI117              bfr                             14           64           176           15          175            177
XI118              bfr                             1            66           45            14          67             173
XI119              bfr                             191          172          163           1           161            166
XI121              bfr                             2            176          169           5           177            36
XI122              bfr                             3            45           35            2           173            44
XI123              bfr                             197          163          32            3           166            42
XI125              bfr                             6            169          28            7           36             37
XI126              bfr                             4            35           174           6           44             34
XI127              bfr                             216          32           164           4           42             165
XI129              bfr                             9            28           170           10          37             162
XI130              bfr                             8            174          178           9           34             167
XI131              bfr                             224          164          178           8           165            162
XI1392             bfr                             323          26           410           259         24             25
XI1393             bfr                             259          412          410           302         20             238
XI1394             bfr                             302          22           304           229         23             50
XI1395             bfr                             229          306          304           230         305            303
XI1396             bfr                             230          313          49            236         48             50
XI1398             bfr                             202          119          206           338         118            205
XI1400             bfr                             204          19           325           273         209            324
XI1401             bfr                             199          325          412           298         324            20
XI1403             bfr                             298          411          22            234         21             23
XI20               bfr                             290          492          494           420         82             493
XI21               bfr                             291          83           78            290         491            79
XI22               bfr                             267          499          54            489         80             52
XI23               bfr                             296          68           322           267         69             55
XI24               bfr                             508          335          438           182         433            130
XI25               bfr                             182          335          436           525         526            131
XI26               bfr                             525          299          434           185         529            132
XI28               bfr                             342          380          126           312         530            127
XI29               bfr                             340          135          128           342         527            443
XI30               bfr                             214          135          134           340         531            427
XI31               bfr                             343          16           124           214         528            125
XI32               bfr                             347          110          462           321         108            109
XI33               bfr                             348          465          107           347         106            463
XI34               bfr                             349          105          104           348         467            466
XI35               bfr                             521          103          102           349         469            468
XI36               bfr                             352          94           483           355         93             482
XI37               bfr                             351          99           98            352         479            478
XI38               bfr                             353          97           480           351         95             96
XI39               bfr                             181          484          91            353         90             92
XI40               bfr                             430          496          502           337         495            75
XI41               bfr                             346          498          503           430         81             73
XI42               bfr                             345          120          454           346         455            453
XI43               bfr                             520          88           86            345         85             87
XI44               bfr                             358          126          110           311         127            108
XI45               bfr                             362          128          465           358         443            106
XI46               bfr                             367          134          105           362         427            467
XI47               bfr                             373          124          103           367         125            469
XI48               bfr                             378          462          94            320         109            93
XI488              bfr                             240          327          242           187         43             241
XI49               bfr                             379          107          99            378         463            479
XI490              bfr                             244          242          40            213         241            41
XI50               bfr                             381          104          97            379         466            95
XI51               bfr                             388          102          484           381         468            90
XI52               bfr                             392          483          496           393         482            495
XI53               bfr                             395          98           498           392         478            81
XI54               bfr                             398          480          120           395         96             455
XI55               bfr                             402          91           88            398         92             85
XI56               bfr                             405          502          501           336         75             76
XI57               bfr                             408          503          501           405         73             74
XI58               bfr                             409          454          71            408         453            76
XI59               bfr                             357          86           71            409         87             74
XI603              bfr                             287          488          83            270         89             491
XI604              bfr                             270          84           492           522         490            82
XI672              bfr                             254          339          256           250         341            255
XI673              bfr                             261          256          31            215         255            262
XI674              bfr                             250          339          441           226         33             435
XI675              bfr                             272          289          29            279         288            30
XI676              bfr                             417          29           461           280         30             457
XI677              bfr                             415          294          27            281         293            407
XI686              bfr                             297          27           333           237         407            332
XI687              bfr                             301          148          411           248         282            21
XI690              bfr                             248          330          143           249         329            309
XI693              bfr                             226          184          488           227         341            89
XI697              bfr                             281          322          308           274         55             56
XI698              bfr                             280          500          506           276         77             505
XI699              bfr                             279          78           500           277         79             77
XI700              bfr                             237          308          46            239         56             47
XI706              bfr                             249          40           307           515         41             51
XI708              bfr                             231          307          233           193         51             232
XI709              bfr                             227          184          84            517         133            490
XI713              bfr                             274          54           264           200         52             53
XI714              bfr                             276          504          70            183         72             509
XI715              bfr                             277          494          504           188         493            72
XI716              bfr                             239          264          327           211         53             43
XI864              bfr                             515          111          146           217         112            144
XI869              bfr                             517          432          519           513         433            518
XI893              bfr                             200          497          121           198         510            122
XI894              bfr                             183          426          450           422         136            444
XI895              bfr                             188          17           426           192         511            136
XI935              bfr                             211          121          115           208         122            460
XI974              bfr                             235          233          313           201         232            48
XI978              bfr                             275          70           499           464         509            80
XI979              bfr                             292          506          68            275         505            69
XI99               bfr                             328          31           385           265         262            383
XI1218             const0                          100          485          223           101         150
XI1376             maj3_KSA_GP_ene_opt             260          310          312           530         527            160                    382        311   142       380       159        158
XI1377             maj3_KSA_GP_ene_opt             316          319          321           160         382            157                    404        320   159       158       403        406
XI1382             maj3_KSA_GP_ene_opt             331          334          355           157         404            155                    419        393   403       406       156        421
XI1383             maj3_KSA_GP_ene_opt             326          323          337           155         419            238                    25         336   156       421       225        225
XI1384             maj3_KSA_sum_ene_opt_boost      514          132          131           130         442            153                    439        189   486       434       436        438        152        440        154        191
XI1385             maj3_KSA_sum_ene_opt_boost      437          442          153           439         451            448                    446        196   195       152       440        154        449        447        445        197
XI1390             maj3_KSA_sum_ene_opt_boost      210          451          448           446         476            474                    472        338   149       449       447        445        475        473        471        216
XI1391             maj3_KSA_sum_ene_opt_boost      207          476          474           472         487            150                    487        219   223       475       473        471        151        151        485        224
XI428              maj_bbb                         263          265          215           251         441            287                    253        435
XI429              maj_bbb                         384          285          295           283         461            292                    284        457
XI438              maj_bbb                         273          246          247           148         333            243                    282        332
XI1088             or_bb                           387          512          429           129         508            431                    371
XI1091             or_bb                           390          481          428           300         486            425                    18
XSUM0              sink                            10           38           170           39          167
XSUM1              sink                            7            171          38            168         39
XSUM2              sink                            5            58           171           59          168
XSUM3              sink                            15           61           58            57          59
XSUM4              sink                            13           0            61            0           57
XI100              spl2                            269          385          140           271         383            386                    272
XI101              spl2                            268          140          391           417         386            389                    295
XI103              spl2                            331          138          139           245         400            401                    252
XI104              spl2                            245          399          397           297         394            396                    247
XI107              spl2                            266          414          418           246         413            416                    286
XI108              spl2                            334          139          194           266         401            137                    507
XI1397             spl2                            201          146          147           202         144            145                    203
XI1399             spl2                            326          194          26            204         137            24                     199
XI1402             spl2                            234          143          306           231         309            305                    235
XI489              spl2                            243          46           330           240         47             329                    244
XI629              spl2                            356          318          399           228         317            394                    415
XI630              spl2                            354          315          318           278         314            317                    285
XI631              spl2                            319          141          138           354         368            400                    356
XI671              spl2                            260          142          258           254         33             257                    261
XI97               spl2                            310          258          350           328         257            344                    269
XI98               spl2                            316          350          141           268         344            368                    370
*end of top cell   maj3_4_bit_KSA_ene_opt_booster


.tran              {{t_step}}ps                    {{end}}ps    {{begin}}ps  {{t_step}}ps
.FiLE              {{out_file_name}}
.print             i(Rac1)
*vac1_tot
.print             nodev                           528          0

.print             i(Rac2)
*vac2_tot
.print             nodev                           531          0

*vac1_DUT
.print             nodev                           527          526
*vac2_DUT
.print             nodev                           530          529