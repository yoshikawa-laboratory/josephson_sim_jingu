.model             jjmod              jj(Rtype=1,  Vg=2.8mV,    Cap=0.064pF,       R0=100ohm,  Rn=17ohm,      Icrit=0.1mA)


.subckt            branch3            1            2            3                  4
*inst name         cell_name          a            b            c                  d
Lip                7                  4            0.312pH
Lp1                1                  6            11.8pH
Lp2                2                  7            10.2pH
Lp3                3                  5            11.8pH
R0                 6                  7            1e-12ohm
R1                 5                  7            1e-12ohm
.ends


.subckt            const0             1            2            11                 12          13
*inst name         cell_name          din          dout         q                  xin         xout
B1                 8                  0            jjmod        area=0.5
B2                 4                  0            jjmod        area=0.5
Kd1                Ld                 L1           -0.128
Kd2                Ld                 L2           -0.135
Kdout              Ld                 Lout         -0.000253
Kdq                Ld                 Lq           -0.00468
Kout               Lq                 Lout         -0.495
Kx1                Lx                 L1           -0.185
Kx2                Lx                 L2           -0.189
Kxd                Lx                 Ld           0.193
Kxout              Lx                 Lout         -7.94e-05
Kxq                Lx                 Lq           -0.00421
L1                 7                  8            1.56pH
L2                 4                  7            1.66pH
Ld                 1                  2            7.49pH
Lout               5                  11           31.2pH
Lq                 7                  0            7.82pH
Lx                 12                 13           7.47pH
R1                 5                  0            1e-12ohm
.ends


.subckt            bfr                1            2            3                  12          13             14
*inst name         cell_name          a            din          dout               q           xin            xout
B1                 9                  0            jjmod        area=0.5
B2                 5                  0            jjmod        area=0.5
Kd1                Ld                 L1           -0.133
Kd2                Ld                 L2           -0.133
Kdout              Ld                 Lout         0.0
Kdq                Ld                 Lq           0.0
Kout               Lq                 Lout         -0.495
Kx1                Lx                 L1           -0.186
Kx2                Lx                 L2           -0.186
Kxd                Lx                 Ld           0.19
Kxout              Lx                 Lout         0.0
Kxq                Lx                 Lq           0.0
L1                 8                  9            1.59pH
L2                 5                  8            1.59pH
Ld                 2                  3            7.45pH
Lin                1                  8            1.23pH
Lout               6                  12           31.2pH
Lq                 8                  0            7.92pH
Lx                 13                 14           7.4pH
R1                 6                  0            1e-12ohm
.ends


.subckt            and_bb             1            2            3                  4           12             13                     14
*inst name         cell_name          a            b            din                dout        q              xin                    xout
XI0                bfr                1            3            8                  9           13             5
XI2                bfr                2            11           4                  10          7              14
XI3                branch3            9            6            10                 12
XI1                const0             8            11           6                  5           7
.ends


.subckt            bias_pair_10um     1            2            3                  4
*inst name         cell_name          a            b            c                  d
*C0                 2                  0            0.00145pF
*C6                 4                  0            0.00144pF
L0                 1                  2            3.46pH
L1                 3                  4            3.73pH
.ends


.subckt            branch2            1            2            3
*inst name         cell_name          a            b            c
Lip                6                  3            0.282pH
Lp1                1                  5            11.0pH
Lp2                2                  4            11.0pH
R0                 5                  6            1e-12ohm
R1                 4                  6            1e-12ohm
.ends


.subckt            spl2               1            2            3                  9           10             11                     12
*inst name         cell_name          a            din          dout               x           xin            xout                   y
XI0                bfr                1            4            6                  7           8              5
XI14               bias_pair_10um     10           8            2                  4
XI15               bias_pair_10um     5            11           6                  3
XI1                branch2            9            12           7
.ends


.subckt            inv                1            2            3                  12          13             14
*inst name         cell_name          a            din          dout               q           xin            xout
B1                 9                  0            jjmod        area=0.6
B2                 5                  0            jjmod        area=0.6
Kd1                Ld                 L1           -0.133
Kd2                Ld                 L2           -0.133
Kdout              Ld                 Lout         0.0
Kdq                Ld                 Lq           0.0
Kout               Lq                 Lout         0.432
Kx1                Lx                 L1           -0.186
Kx2                Lx                 L2           -0.186
Kxd                Lx                 Ld           0.19
Kxout              Lx                 Lout         0.0
Kxq                Lx                 Lq           0.0
L1                 8                  9            1.59pH
L2                 5                  8            1.59pH
Ld                 2                  3            7.44pH
Lin                1                  8            1.24pH
Lout               6                  12           31.0pH
Lq                 8                  0            6.49pH
Lx                 13                 14           7.39pH
R1                 6                  0            1e-12ohm
.ends


.subckt            maj_bbi            1            2            3                  4           5              13                     14    15
*inst name         cell_name          a            b            c                  din         dout           q                      xin   xout
XI0                bfr                1            4            9                  11          14             6
XI1                bfr                2            9            12                 7           6              8
XI3                branch3            11           7            10                 13
XI2                inv                3            12           5                  10          8              15
.ends


.subckt            bias_pair_20um     1            2            3                  4
*inst name         cell_name          a            b            c                  d
XI0                bias_pair_10um     1            6            3                  5
XI1                bias_pair_10um     6            2            5                  4
.ends


.subckt            bfrL               1            2            3                  12          13             14
*inst name         cell_name          a            din          dout               q           xin            xout
B1                 9                  0            jjmod        area=1.0
B2                 5                  0            jjmod        area=1.0
Kd1                Ld                 L1           -0.135
Kd2                Ld                 L2           -0.135
Kdout              Ld                 Lout         0.0
Kdq                Ld                 Lq           0.0
Kout               Lq                 Lout         -0.495
Kx1                Lx                 L1           -0.187
Kx2                Lx                 L2           -0.187
Kxd                Lx                 Ld           0.192
Kxout              Lx                 Lout         0.0
Kxq                Lx                 Lq           0.0
L1                 8                  9            1.59pH
L2                 5                  8            1.59pH
Ld                 2                  3            7.43pH
Lin                1                  8            1.24pH
Lout               6                  12           31.1pH
Lq                 8                  0            7.92pH
Lx                 13                 14           7.38pH
R1                 6                  0            1e-12ohm
.ends


.subckt            spl3L              1            2            3                  9           10             11                     12    13
*inst name         cell_name          a            din          dout               x           xin            xout                   y     z
XI0                bfrL               1            4            6                  7           8              5
XI14               bias_pair_20um     10           8            2                  4
XI15               bias_pair_20um     5            11           6                  3
XI1                branch3            9            12           13                 7
.ends


.subckt            maj_bib            1            2            3                  4           5              13                     14    15
*inst name         cell_name          a            b            c                  din         dout           q                      xin   xout
XI0                bfr                1            4            9                  11          14             6
XI2                bfr                3            7            5                  10          8              15
XI3                branch3            11           12           10                 13
XI1                inv                2            9            7                  12          6              8
.ends


.subckt            maj_ibb            1            2            3                  4           5              13                     14    15
*inst name         cell_name          a            b            c                  din         dout           q                      xin   xout
XI1                bfr                2            8            10                 12          6              7
XI2                bfr                3            10           5                  9           7              15
XI3                branch3            11           12           9                  13
XI0                inv                1            4            8                  11          14             6
.ends


.subckt            maj_bbb            1            2            3                  4           5              13                     14    15
*inst name         cell_name          a            b            c                  din         dout           q                      xin   xout
XI0                bfr                1            4            8                  11          14             6
XI1                bfr                2            8            10                 12          6              7
XI2                bfr                3            10           5                  9           7              15
XI3                branch3            11           12           9                  13
.ends


.subckt            sink               1            2            3                  10          11
*inst name         cell_name          a            din          dout               xin         xout
B1                 8                  0            jjmod        area=0.5
B2                 5                  0            jjmod        area=0.5
Kd1                Ld                 L1           -0.133
Kd2                Ld                 L2           -0.133
Kdq                Ld                 Lq           0.0
Kx1                Lx                 L1           -0.186
Kx2                Lx                 L2           -0.186
Kxd                Lx                 Ld           0.19
Kxq                Lx                 Lq           0.0
L1                 7                  8            1.59pH
L2                 5                  7            1.59pH
Ld                 2                  3            7.45pH
Lin                1                  7            1.23pH
Lq                 7                  0            7.92pH
Lx                 10                 11           7.4pH
.ends


.subckt            and_bi             1            2            3                  4           12             13                     14
*inst name         cell_name          a            b            din                dout        q              xin                    xout
XI0                bfr                1            3            8                  9           13             5
XI3                branch3            9            7            10                 12
XI1                const0             8            11           7                  5           6
XI2                inv                2            11           4                  10          6              14
.ends


.subckt            const1             1            2            7                  8           9
*inst name         cell_name          din          dout         q                  xin         xout
L1                 8                  4            0.01pH
L2                 6                  9            0.01pH
L3                 1                  3            0.01pH
L4                 5                  2            0.01pH
XI0                const0             5            3            7                  6           4
.ends


.subckt            or_bb              1            2            3                  4           12             13                     14
*inst name         cell_name          a            b            din                dout        q              xin                    xout
XI0                bfr                1            3            8                  9           13             5
XI2                bfr                2            11           4                  10          6              14
XI3                branch3            9            7            10                 12
XI1                const1             8            11           7                  5           6
.ends


*this is top cell  16bit_RCA_ene_opt
R37                3186               2134         1000.0ohm
R38                3210               3428         1000.0ohm
R39                2277               3417         1000.0ohm
R40                3255               375          1000.0ohm
R41                526                1596         1000.0ohm
R42                1567               707          1000.0ohm
R43                596                1467         1000.0ohm
R44                288                252          1000.0ohm
R45                276                254          1000.0ohm
R46                2933               3074         1000.0ohm
R47                3028               237          1000.0ohm
R48                272                239          1000.0ohm
R49                268                238          1000.0ohm
R50                2760               251          1000.0ohm
R51                264                3199         1000.0ohm
R52                3267               3295         1000.0ohm
R53                3145               2161         1000.0ohm
R54                3244               3444         1000.0ohm
R55                2228               3440         1000.0ohm
R56                747                629          1000.0ohm
R57                765                678          1000.0ohm
R58                1491               1483         1000.0ohm
R59                1454               1518         1000.0ohm
R60                286                256          1000.0ohm
R61                274                2618         1000.0ohm
R62                281                2896         1000.0ohm
R63                3204               236          1000.0ohm
R64                270                2794         1000.0ohm
R65                266                247          1000.0ohm
R66                260                249          1000.0ohm
R67                262                230          1000.0ohm
R68                400                1824         1000.0ohm
Rac1               3236               3497         100000.0ohm
Rac2               3054               3500         100000.0ohm
Rdc1               3273               947          100000.0ohm
V10                3255               0            PWL          (0ps 0mV 20ps {{input[0]}})
V11                747                0            PWL          (0ps 0mV 20ps {{input[1]}})
V12                526                0            PWL          (0ps 0mV 20ps {{input[2]}})
V13                765                0            PWL          (0ps 0mV 20ps {{input[3]}})
V14                1567               0            PWL          (0ps 0mV 20ps {{input[4]}})
V15                1491               0            PWL          (0ps 0mV 20ps {{input[5]}})
V16                596                0            PWL          (0ps 0mV 20ps {{input[6]}})
V17                1454               0            PWL          (0ps 0mV 20ps {{input[7]}})
V19                400                0            PWL          (0ps 0mV 20ps {{input[8]}})
V21                288                0            PWL          (0ps 0mV 20ps {{input[9]}})
V22                286                0            PWL          (0ps 0mV 20ps {{input[10]}})
V23                276                0            PWL          (0ps 0mV 20ps {{input[11]}})
V24                274                0            PWL          (0ps 0mV 20ps {{input[12]}})
V25                2933               0            PWL          (0ps 0mV 20ps {{input[13]}})
V26                281                0            PWL          (0ps 0mV 20ps {{input[14]}})
V27                3028               0            PWL          (0ps 0mV 20ps {{input[15]}})
V28                3204               0            PWL          (0ps 0mV 20ps {{input[16]}})
V29                272                0            PWL          (0ps 0mV 20ps {{input[17]}})
V3                 3267               0            PWL          (0ps 0mV 20ps {{input[18]}})
V30                270                0            PWL          (0ps 0mV 20ps {{input[19]}})
V31                268                0            PWL          (0ps 0mV 20ps {{input[20]}})
V32                266                0            PWL          (0ps 0mV 20ps {{input[21]}})
V33                2760               0            PWL          (0ps 0mV 20ps {{input[22]}})
V34                260                0            PWL          (0ps 0mV 20ps {{input[23]}})
V35                264                0            PWL          (0ps 0mV 20ps {{input[24]}})
V36                262                0            PWL          (0ps 0mV 20ps {{input[25]}})
V4                 3186               0            PWL          (0ps 0mV 20ps {{input[26]}})
V5                 3145               0            PWL          (0ps 0mV 20ps {{input[27]}})
V6                 3210               0            PWL          (0ps 0mV 20ps {{input[28]}})
V7                 3244               0            PWL          (0ps 0mV 20ps {{input[29]}})
V8                 2277               0            PWL          (0ps 0mV 20ps {{input[30]}})
V9                 2228               0            PWL          (0ps 0mV 20ps {{input[31]}})
VDC                3273               0            PWL          (0ps               0mV         20ps           113000mV)
VAC1               3236               0            SIN          (0                 81000mV     {{freq}}MEGHz  {{40+period|int/4}}ps  0)
VAC2               3054               0            SIN          (0                 81000mV     {{freq}}MEGHz  40ps                   0)
XI0                and_bb             1930         2640         2093               481         2284           2031                   869
XI1201             and_bi             2143         2225         687                2292        2229           1135                   2095
XI156              and_bi             1994         3445         2292               2111        2179           2095                   3275
XI100              bfr                3344         2454         2425               3439        427            2386
XI1000             bfr                256          916          911                231         917            912
XI1001             bfr                632          909          907                150         891            908
XI1002             bfr                529          907          906                3016        908            903
XI1003             bfr                716          906          904                3069        903            901
XI1004             bfr                517          904          902                2899        901            898
XI1005             bfr                1            902          900                107         898            896
XI1006             bfr                708          900          897                2676        896            894
XI1007             bfr                682          897          876                2844        894            895
XI1008             bfr                775          3147         909                2981        395            891
XI1009             bfr                150          890          888                2943        887            889
XI101              bfr                87           2455         2454               643         355            427
XI1010             bfr                2899         886          885                3167        883            878
XI1011             bfr                3069         881          886                3085        882            883
XI1012             bfr                3016         888          881                3035        889            882
XI1013             bfr                107          885          875                2777        878            879
XI1014             bfr                2844         877          876                2719        874            3443
XI1015             bfr                2676         875          877                2502        879            874
XI1016             bfr                2981         442          890                2680        872            887
XI1017             bfr                2680         871          870                2843        1687           860
XI1018             bfr                3035         861          867                2948        866            868
XI1019             bfr                3085         867          865                3106        868            862
XI102              bfr                3421         3452         2455               3426        354            355
XI1020             bfr                3167         865          856                53          862            864
XI1021             bfr                2943         870          861                3059        860            866
XI1022             bfr                2502         854          859                2764        855            857
XI1023             bfr                2719         859          833                2613        857            818
XI1024             bfr                2777         856          854                47          864            855
XI1025             bfr                2843         853          851                2520        849            852
XI1026             bfr                2948         840          847                3110        841            848
XI1027             bfr                3106         847          845                2683        848            846
XI1028             bfr                53           845          842                17          846            843
XI1029             bfr                3059         851          840                2552        852            841
XI103              bfr                3356         441          2434               115         2426           421
XI1030             bfr                2764         839          837                3046        835            838
XI1031             bfr                2613         837          833                8           838            834
XI1032             bfr                47           842          839                2867        843            835
XI1033             bfr                2520         1846         830                3003        1847           822
XI1034             bfr                3110         823          829                3480        824            826
XI1035             bfr                2683         829          825                3209        826            828
XI1036             bfr                17           825          816                2643        828            813
XI1037             bfr                2552         830          823                2755        822            824
XI1038             bfr                3046         821          819                2690        815            817
XI1039             bfr                8            819          796                2830        817            818
XI104              bfr                3429         2428         441                301         430            2426
XI1040             bfr                2867         816          821                2756        813            815
XI1041             bfr                3003         812          811                2737        810            800
XI1042             bfr                3480         801          808                3450        807            809
XI1043             bfr                3209         808          805                2686        809            802
XI1044             bfr                2643         805          803                2984        802            804
XI1045             bfr                2755         811          801                3200        800            807
XI1046             bfr                2690         799          797                3432        794            798
XI1047             bfr                2830         797          796                2572        798            834
XI1048             bfr                2756         803          799                2931        804            794
XI1049             bfr                2737         793          2721               2770        1843           792
XI105              bfr                3337         353          2428               3375        2443           430
XI1050             bfr                3450         2841         3014               3404        2784           2723
XI1051             bfr                2686         3014         785                2926        2723           2722
XI1052             bfr                2984         785          3060               2670        2722           770
XI1053             bfr                3200         2721         2841               3182        792            2784
XI1054             bfr                3432         2780         776                2923        2634           2588
XI1055             bfr                2572         776          2887               3133        2588           2968
XI1056             bfr                2931         3060         2780               2940        770            2634
XI1057             bfr                2770         1848         2936               2667        1849           751
XI1058             bfr                3404         2576         2945               2635        2878           2837
XI1059             bfr                2926         2945         3038               2506        2837           2658
XI106              bfr                235          458          353                3344        2442           2443
XI1060             bfr                2670         3038         2865               3324        2658           757
XI1061             bfr                3182         2936         2576               2656        751            2878
XI1062             bfr                2923         750          3135               2507        2565           2982
XI1063             bfr                3133         3135         2887               2942        2982           2869
XI1064             bfr                2940         2865         750                2557        757            2565
XI1065             bfr                2667         1836         731                2939        1837           740
XI1066             bfr                2635         3030         2759               2495        2740           3045
XI1067             bfr                2506         2759         2515               3052        3045           2688
XI1068             bfr                3324         2515         733                2853        2688           734
XI1069             bfr                2656         731          3030               3075        740            2740
XI107              bfr                3446         3361         458                87          3390           2442
XI1070             bfr                2507         3032         726                2697        2806           2804
XI1071             bfr                2942         726          693                2849        2804           2968
XI1072             bfr                2557         733          3032               3154        734            2806
XI1073             bfr                2939         1838         2593               2960        1839           2501
XI1074             bfr                2495         2993         2578               2532        3124           712
XI1075             bfr                3052         2578         2742               2665        712            2753
XI1076             bfr                2853         2742         2928               3109        2753           3192
XI1077             bfr                3075         2593         2993               2819        2501           3124
XI1078             bfr                2697         699          3048               3012        696            692
XI1079             bfr                2849         3048         693                2415        692            2869
XI108              bfr                3433         424          3361               3421        2422           3390
XI1080             bfr                3154         2928         699                3019        3192           696
XI1081             bfr                2960         1998         2765               2674        2725           3123
XI1082             bfr                2532         672          2796               2566        2696           2707
XI1083             bfr                2665         2796         2814               2523        2707           679
XI1084             bfr                3109         2814         675                2493        679            660
XI1085             bfr                2819         2765         672                2791        3123           2696
XI1086             bfr                3012         2546         2644               3207        667            2510
XI1087             bfr                2415         2644         664                3100        2510           2575
XI1088             bfr                3019         675          2546               2808        660            667
XI1089             bfr                2674         2000         658                2795        2001           649
XI109              bfr                3335         2398         3438               62          357            376
XI1090             bfr                2566         3092         656                1977        2662           657
XI1091             bfr                2523         656          3174               2861        657            2592
XI1092             bfr                2493         3174         653                1862        2592           2561
XI1093             bfr                2791         658          3092               3129        649            2662
XI1094             bfr                3207         2763         647                2965        2994           3063
XI1095             bfr                3100         647          664                2716        3063           2836
XI1096             bfr                2808         653          2763               2583        2561           2994
XI1097             bfr                2795         2903         2959               2620        1995           2847
XI1098             bfr                1977         623          2980               2852        2851           2499
XI1099             bfr                2861         2980         2642               3094        2499           2601
XI110              bfr                273          358          2398               78          463            357
XI1100             bfr                1862         2642         628                2559        2601           2781
XI1101             bfr                3129         2959         623                2992        2847           2851
XI1102             bfr                2965         2659         3070               2585        619            616
XI1103             bfr                2716         3070         2652               3183        616            2575
XI1104             bfr                2583         628          2659               2886        2781           619
XI1105             bfr                2620         1992         612                2607        1993           613
XI1106             bfr                2852         2714         609                2617        2700           606
XI1107             bfr                3094         609          3018               2998        606            2788
XI1108             bfr                2559         3018         2741               2769        2788           3082
XI1109             bfr                2992         612          2714               2685        613            2700
XI111              bfr                283          2436         358                1088        2437           463
XI1110             bfr                2585         589          593                2505        594            591
XI1111             bfr                3183         593          2652               2639        591            2836
XI1112             bfr                2886         2741         589                3128        3082           594
XI1113             bfr                2607         587          584                2543        2537           3036
XI1114             bfr                2617         3166         3058               2612        2990           2967
XI1115             bfr                2998         3058         3095               2535        2967           2542
XI1116             bfr                2769         3095         574                2531        2542           2738
XI1117             bfr                2685         584          3166               2630        3036           2990
XI1118             bfr                2505         571          567                3049        568            2678
XI1119             bfr                2639         567          541                2811        2678           3495
XI112              bfr                3439         2438         2436               20          443            2437
XI1120             bfr                3128         574          571                2888        2738           568
XI1121             bfr                2543         563          2649               2875        3000           2827
XI1122             bfr                2612         559          2577               2           2962           3157
XI1123             bfr                2535         2577         2545               2560        3157           550
XI1124             bfr                2531         2545         539                3040        550            535
XI1125             bfr                2630         2649         559                2771        2827           2962
XI1126             bfr                3049         2606         543                2975        537            2704
XI1127             bfr                2811         543          541                3107        2704           3498
XI1128             bfr                2888         539          2606               3008        535            537
XI113              bfr                643          3422         2438               132         3317           443
XI1137             bfr                258          2631         2136               257         488            502
XI1138             bfr                259          2631         3050               258         3105           2138
XI114              bfr                3426         471          3422               245         3457           3317
XI1140             bfr                2664         496          2720               2490        468            495
XI1141             bfr                2540         469          2774               2664        2874           435
XI1142             bfr                2490         496          2137               259         488            2987
XI1159             bfr                3411         3379         3241               3299        3280           3300
XI1160             bfr                3299         3408         3367               3401        3396           3261
XI1162             bfr                3364         3367         3388               3333        3261           3312
XI1163             bfr                25           3241         3398               3364        3300           3362
XI1165             bfr                3399         3388         3265               33          3312           3389
XI1166             bfr                3320         3398         3381               3399        3362           3260
XI1168             bfr                32           3265         3410               3340        3389           3341
XI1169             bfr                3372         3381         3412               32          3260           3363
XI117              bfr                3490         3276         2400               1252        2450           2399
XI1171             bfr                3357         3412         3371               30          3363           3394
XI1172             bfr                30           3410         3403               31          3341           3332
XI1174             bfr                28           3371         2812               3407        3394           3298
XI1175             bfr                3407         3403         3348               3383        3332           3354
XI1177             bfr                3246         2812         504                34          3298           3498
XI1178             bfr                34           3348         3291               22          3354           0
XI118              bfr                1252         483          391                2766        2453           2408
XI1183             bfr                23           2012         3408               3228        2991           3396
XI1184             bfr                3339         531          3379               23          3250           3280
XI1186             bfr                2875         2007         3413               3339        2008           3229
XI1187             bfr                2771         3413         3352               3411        3229           3377
XI1188             bfr                2            3352         521                25          3377           524
XI1189             bfr                2560         521          516                3320        524            515
XI119              bfr                3302         2400         2988               2911        2399           3358
XI1190             bfr                3040         516          3308               3372        515            510
XI1191             bfr                3008         3308         3326               3357        510            512
XI1192             bfr                2975         3326         506                28          512            3345
XI1193             bfr                3107         506          504                3246        3345           3495
XI120              bfr                1861         482          2872               3302        383            385
XI121              bfr                2911         391          3287               3314        2408           2409
XI122              bfr                3493         3349         1109               1861        392            2414
XI123              bfr                3449         2988         405                3385        3358           3435
XI124              bfr                3385         3287         405                3420        2409           2189
XI125              bfr                141          1109         2439               44          2414           3455
XI126              bfr                3494         2458         2892               77          2457           3455
XI127              bfr                44           2872         2439               3449        385            2901
XI128              bfr                77           407          2892               141         479            2901
XI129              bfr                20           26           2446               363         2913           2444
XI130              bfr                1088         2446         2445               411         2444           2405
XI131              bfr                62           387          2417               225         2406           2418
XI132              bfr                78           2445         387                307         2405           2406
XI133              bfr                831          390          291                953         2407           263
XI134              bfr                132          2435         26                 831         394            2913
XI135              bfr                411          448          2413               522         449            2411
XI136              bfr                522          326          379                680         2424           198
XI137              bfr                245          255          2435               763         46             394
XI138              bfr                307          2413         2394               3491        2411           401
XI139              bfr                225          2394         481                3492        401            869
XI140              bfr                680          2391         2388               3489        2387           486
XI141              bfr                603          3281         2391               3488        2383           2387
XI142              bfr                1253         498          3272               3485        84             380
XI143              bfr                1312         3272         485                3486        380            3346
XI144              bfr                1134         2287         436                1253        368            434
XI145              bfr                1194         436          2174               1312        434            2429
XI146              bfr                1015         2461         2404               1134        2459           2403
XI147              bfr                892          2433         413                1015        29             2432
XI148              bfr                953          413          370                1074        2432           373
XI149              bfr                1074         2404         3281               1194        2403           2383
XI150              bfr                464          370          326                603         373            2424
XI151              bfr                763          36           390                892         2401           2407
XI152              bfr                363          291          448                464         263            449
XI168              bfr                554          284          2375               570         3269           2376
XI169              bfr                570          2373         278                632         2372           2368
XI175              bfr                530          2375         2371               507         2376           2366
XI176              bfr                544          261          2364               530         2369           2363
XI177              bfr                507          278          2365               529         2368           234
XI182              bfr                665          2371         3400               569         2366           2169
XI183              bfr                569          2365         3395               716         234            3391
XI184              bfr                484          2364         3351               665         2363           233
XI186              bfr                685          223          210                475         1534           207
XI187              bfr                475          1573         2357               478         2360           215
XI188              bfr                552          2359         221                685         1494           222
XI190              bfr                460          2357         476                455         215            3330
XI191              bfr                778          221          2355               447         222            213
XI192              bfr                447          210          369                460         207            209
XI194              bfr                425          2355         2354               433         213            2352
XI200              bfr                669          2354         3329               788         2352           3328
XI212              bfr                702          404          199                544         566            2350
XI220              bfr                167          199          2351               484         2350           2154
XI221              bfr                780          2349         2347               167         3327           2168
XI222              bfr                160          191          2167               780         525            756
XI226              bfr                124          2346         2345               575         2344           178
XI227              bfr                575          185          2340               552         1455           170
XI228              bfr                3            1378         182                124         1379           2341
XI229              bfr                599          2345         2342               540         178            180
XI230              bfr                646          182          2338               599         2341           2337
XI231              bfr                540          2340         171                778         170            166
XI232              bfr                99           171          168                425         166            2332
XI233              bfr                3471         2338         164                94          2337           149
XI234              bfr                94           2342         161                99          180            2334
XI235              bfr                85           161          2335               545         2334           2326
XI236              bfr                545          168          728                669         2332           156
XI237              bfr                3466         164          2331               85          149            147
XI238              bfr                761          2331         2330               700         147            2324
XI239              bfr                700          2335         145                82          2326           138
XI240              bfr                74           145          686                71          138            140
XI241              bfr                752          2330         136                74          2324           3213
XI249              bfr                3482         183          2323               3           1337           2321
XI250              bfr                556          1298         129                3482        181            130
XI251              bfr                3475         2323         2319               646         2321           2318
XI252              bfr                695          129          122                3475        130            118
XI253              bfr                3386         122          2320               3468        118            109
XI254              bfr                3468         2319         2317               3471        2318           113
XI255              bfr                3462         2317         2315               3466        113            2313
XI256              bfr                3368         2320         110                3462        109            111
XI257              bfr                694          110          106                3451        111            2310
XI258              bfr                3451         2315         2312               761         2313           2311
XI259              bfr                676          2312         2308               752         2311           93
XI260              bfr                3336         106          92                 676         2310           89
XI261              bfr                742          96           3365               3424        95             487
XI262              bfr                3437         2308         96                 3442        93             95
XI263              bfr                721          92           90                 3437        89             91
XI264              bfr                640          90           393                742         91             88
XI265              bfr                3415         2306         86                 556         1261           76
XI266              bfr                3303         2305         2302               721         2301           2303
XI267              bfr                620          2302         498                640         2303           84
XI268              bfr                3338         83           2305               3336        2299           2301
XI269              bfr                3343         2297         83                 694         81             2299
XI270              bfr                648          2298         2297               3368        2294           81
XI271              bfr                720          79           2298               3386        2293           2294
XI272              bfr                715          86           79                 695         76             2293
XI273              bfr                644          2291         2289               3303        75             2290
XI274              bfr                2102         2289         2287               620         2290           368
XI275              bfr                3277         1223         2285               3415        2286           73
XI276              bfr                3253         2285         72                 715         73             70
XI277              bfr                3231         72           69                 720         70             2281
XI278              bfr                3072         69           2280               648         2281           66
XI279              bfr                2912         2280         68                 3343        66             2279
XI280              bfr                2681         68           2291               3338        2279           75
XI281              bfr                719          2278         2267               3277        2275           2265
XI282              bfr                626          2274         64                 644         63             2272
XI283              bfr                2041         64           2461               2102        2272           2459
XI284              bfr                579          60           2274               2681        61             63
XI285              bfr                754          2269         60                 2912        2271           61
XI286              bfr                565          2270         2269               3072        2268           2271
XI287              bfr                3162         58           2270               3231        59             2268
XI288              bfr                3242         2267         58                 3253        2265           59
XI289              bfr                677          16           2238               626         56             27
XI290              bfr                578          2264         2254               759         54             55
XI291              bfr                558          51           2264               2218        52             54
XI292              bfr                577          2262         51                 2295        49             52
XI293              bfr                500          50           2262               2361        48             49
XI294              bfr                2016         2260         50                 724         2259           48
XI295              bfr                1984         2258         2260               2517        2257           2259
XI296              bfr                501          2253         255                598         43             46
XI297              bfr                661          2254         2253               766         55             43
XI298              bfr                724          42           41                 2451        2251           2250
XI299              bfr                2361         41           39                 2389        2250           40
XI300              bfr                2295         39           38                 2328        40             2248
XI301              bfr                2218         38           2247               2255        2248           2245
XI302              bfr                759          2247         2241               2160        2245           2246
XI303              bfr                598          2244         36                 633         2242           2401
XI304              bfr                766          2241         2244               677         2246           2242
XI305              bfr                2517         2240         42                 2604        2239           2251
XI306              bfr                633          2238         2433               2041        27             29
XI307              bfr                2604         1144         2235               719         24             2236
XI308              bfr                2451         2235         2234               3242        2236           19
XI309              bfr                2389         2234         2232               3162        19             21
XI310              bfr                2328         2232         2230               565         21             2231
XI311              bfr                2255         2230         18                 754         2231           15
XI312              bfr                2160         18           16                 579         15             56
XI313              bfr                781          1029         2222               1984        1030           14
XI314              bfr                1518         913          7                  1991        914            2227
XI315              bfr                1991         951          10                 760         952            2226
XI316              bfr                760          991          2223               781         992            2224
XI317              bfr                652          2223         3484               654         2224           3483
XI318              bfr                654          2222         2217               2016        14             11
XI319              bfr                704          10           2219               652         2226           9
XI320              bfr                1467         7            6                  704         2227           2220
XI321              bfr                2028         2219         4                  605         9              5
XI322              bfr                519          2217         2215               500         11             2216
XI323              bfr                605          3484         2211               519         3483           3478
XI324              bfr                1483         6            3481               2028        2220           2212
XI325              bfr                714          2215         2206               577         2216           2214
XI326              bfr                707          3481         3472               703         2212           2205
XI327              bfr                617          2211         2208               714         3478           3479
XI328              bfr                703          4            3476               617         5              3477
XI329              bfr                622          3476         2203               637         3477           2209
XI330              bfr                637          2208         3474               666         3479           2207
XI331              bfr                666          2206         2202               558         2214           3473
XI332              bfr                678          3472         3467               622         2205           3470
XI333              bfr                1924         3474         3464               546         2207           3461
XI334              bfr                1939         2203         2200               1924        2209           3469
XI335              bfr                1596         3467         3460               1939        3470           3458
XI336              bfr                546          2202         2199               578         3473           2197
XI337              bfr                511          2200         3456               492         3469           3454
XI338              bfr                490          2199         2195               661         2197           3465
XI339              bfr                492          3464         3453               490         3461           3463
XI340              bfr                629          3460         3459               511         3458           2196
XI341              bfr                743          2195         471                501         3465           3457
XI342              bfr                1600         3456         424                1607        3454           2422
XI343              bfr                1607         3453         3452               743         3463           354
XI344              bfr                375          3459         2193               1600        2196           2430
XI359              bfr                499          772          2192               625         3434           895
XI360              bfr                625          3431         2192               682         2183           3443
XI361              bfr                608          3427         573                602         489            729
XI362              bfr                601          3425         573                608         2190           784
XI363              bfr                718          3423         2187               601         3436           2189
XI364              bfr                3420         2188         2187               718         2186           3435
XI365              bfr                736          2185         772                758         3419           3434
XI366              bfr                758          2184         3431               708         3430           2183
XI367              bfr                555          2172         3427               630         2173           489
XI368              bfr                536          2182         3425               555         2181           2190
XI369              bfr                642          2180         3423               536         783            3436
XI370              bfr                3314         2178         2188               642         2176           2186
XI371              bfr                497          2175         2185               503         3397           3419
XI372              bfr                503          771          2184               1           3393           3430
XI373              bfr                592          749          2172               787         650            2173
XI374              bfr                786          655          2182               592         2165           2181
XI375              bfr                2766         2171         2178               745         3405           2176
XI376              bfr                745          3376         2180               786         3378           783
XI377              bfr                576          3400         2175               610         2169           3397
XI378              bfr                610          3395         771                517         3391           3393
XI379              bfr                557          2347         749                549         2168           650
XI380              bfr                590          2167         655                557         756            2165
XI381              bfr                1619         3387         2171               583         3382           3405
XI382              bfr                583          472          3376               590         473            3378
XI383              bfr                602          2163         3374               508         585            784
XI384              bfr                508          2159         3374               499         2162           729
XI385              bfr                630          2158         2163               2327        769            585
XI386              bfr                2327         2155         2159               736         3359           2162
XI387              bfr                787          3366         2158               513         2156           769
XI388              bfr                513          2153         2155               497         3350           3359
XI389              bfr                549          2351         3366               710         2154           2156
XI390              bfr                710          3351         2153               576         233            3350
XI393              bfr                3232         2152         2151               2978        2150           2142
XI394              bfr                2978         2149         2145               2953        2146           2148
XI399              bfr                3159         2145         2144               2950        2148           466
XI400              bfr                2894         2151         346                3159        2142           3142
XI402              bfr                3104         3050         2139               155         2138           2140
XI403              bfr                3313         2137         2133               3104        2987           2130
XI404              bfr                155          2136         2129               154         502            2135
XI417              bfr                2768         2133         2131               2839        2130           2132
XI418              bfr                2689         2129         2128               159         2135           2119
XI419              bfr                2839         2139         2125               2689        2140           2126
XI420              bfr                3288         2921         2124               3290        403            2114
XI421              bfr                3290         467          2109               2768        2121           2123
XI430              bfr                2616         2131         2104               3137        2132           2099
XI431              bfr                2521         2128         2120               165         2119           2096
XI432              bfr                3137         2125         2117               2521        2126           2092
XI433              bfr                3274         2124         2115               2653        2114           2116
XI434              bfr                3198         2113         2112               3274        2110           2087
XI435              bfr                2653         2109         2107               2616        2123           2108
XI436              bfr                2729         2106         2086               3198        2105           2084
XI441              bfr                3259         2104         2100               2947        2099           2101
XI442              bfr                177          2120         2097               176         2096           2098
XI443              bfr                2947         2117         2075               177         2092           2094
XI444              bfr                2695         2115         2091               2666        2116           2068
XI445              bfr                2666         2107         2090               3259        2108           2067
XI446              bfr                2815         2112         2060               2695        2087           2088
XI447              bfr                3262         2086         2085               2815        2084           2061
XI448              bfr                2570         2083         2081               3262        2079           2082
XI449              bfr                2691         2078         2077               2570        2076           2063
XI451              bfr                173          2075         2057               175         2094           2074
XI452              bfr                175          2097         2072               174         2098           2056
XI453              bfr                3252         2100         2055               173         2101           2071
XI454              bfr                3258         2091         2070               3257        2068           2050
XI455              bfr                3257         2090         2049               3252        2067           2048
XI456              bfr                3256         2081         2066               3254        2082           2046
XI457              bfr                3130         2077         2045               3256        2063           2064
XI458              bfr                3254         2085         2062               2929        2061           2039
XI459              bfr                2929         2060         2038               3258        2088           2059
XI461              bfr                2761         2057         2036               3216        2074           2033
XI462              bfr                3216         2072         2032               3044        2056           2029
XI463              bfr                2862         2055         2052               2761        2071           2053
XI464              bfr                3251         2070         2051               3247        2050           2027
XI465              bfr                3247         2049         2026               2862        2048           2024
XI466              bfr                2743         2066         2023               3068        2046           2047
XI467              bfr                3206         2045         2043               2743        2064           2044
XI468              bfr                3068         2062         2040               3248        2039           2018
XI469              bfr                3248         2038         2017               3251        2059           2037
XI471              bfr                2951         2036         2013               3138        2033           2035
XI472              bfr                3138         2032         2030               184         2029           2010
XI473              bfr                3239         2052         2009               2951        2053           2006
XI474              bfr                3245         2051         2005               3152        2027           2004
XI475              bfr                3152         2026         2025               3239        2024           2003
XI476              bfr                3243         2023         2002               2734        2047           1999
XI477              bfr                2598         2043         2021               3243        2044           1996
XI478              bfr                2734         2040         2019               3240        2018           2020
XI479              bfr                3240         2017         2014               3245        2037           2015
XI481              bfr                2574         2013         531                2648        2035           3250
XI482              bfr                2648         2030         2012               3024        2010           2991
XI483              bfr                2669         2009         2007               2574        2006           2008
XI484              bfr                3238         2005         587                3237        2004           2537
XI485              bfr                3237         2025         563                2669        2003           3000
XI486              bfr                2509         2002         2000               3234        1999           2001
XI487              bfr                2358         2021         1998               2509        1996           2725
XI488              bfr                3234         2019         2903               2845        2020           1995
XI489              bfr                2845         2014         1992               3238        2015           1993
XI491              bfr                3151         2152         1974               3232        2146           1990
XI492              bfr                3221         1989         1987               3227        1986           1988
XI493              bfr                3227         1989         1985               3151        2150           1967
XI494              bfr                2935         1983         1970               3221        1981           1982
XI495              bfr                3202         1983         1980               2935        1986           1965
XI496              bfr                3194         1979         1976               3202        1981           1963
XI497              bfr                2909         1979         1962               3194        1975           1961
XI498              bfr                3178         1974         1972               2894        1990           1973
XI499              bfr                3163         1987         1955               3169        1988           1952
XI500              bfr                3153         1970         1956               3163        1982           1969
XI501              bfr                3169         1985         1959               3178        1967           1957
XI502              bfr                2705         1980         1966               3153        1965           1947
XI503              bfr                2611         1976         1951               2705        1963           1949
XI504              bfr                2946         1962         1946               2611        1961           1943
XI505              bfr                3117         1972         1960               3127        1973           1941
XI506              bfr                3108         1959         1937               3117        1957           1935
XI507              bfr                3091         1956         1934               3099        1969           1932
XI508              bfr                3099         1955         1954               3108        1952           1938
XI509              bfr                3073         1951         1950               2904        1949           1927
XI510              bfr                2904         1966         1931               3091        1947           1948
XI511              bfr                2805         1946         1944               3073        1943           1923
XI512              bfr                2498         1960         1942               3064        1941           461
XI513              bfr                2567         1954         1920               2974        1938           1940
XI514              bfr                2974         1937         1936               2498        1935           2679
XI515              bfr                3208         1934         1933               2567        1932           1921
XI516              bfr                3195         1931         1915               3208        1948           1914
XI517              bfr                3013         1950         1928               3195        1927           1929
XI518              bfr                2288         1944         1925               3013        1923           1926
XI519              bfr                2979         1933         1908               2989        1921           1922
XI520              bfr                2989         1920         1911               3103        1940           1909
XI521              bfr                2651         1928         1916               3113        1929           1917
XI522              bfr                3113         1915         1907               2979        1914           1905
XI523              bfr                2868         1925         1913               2651        1926           1902
XI527              bfr                2907         1911         1910               2731        1909           2881
XI528              bfr                2672         1908         331                2907        1922           3180
XI529              bfr                2587         1907         1901               2672        1905           1898
XI530              bfr                3188         1916         1897               2587        1917           1896
XI531              bfr                2823         1913         1903               3188        1902           1904
XI534              bfr                2772         1901         1899               2813        1898           1900
XI535              bfr                2938         1897         1893               2772        1896           1890
XI536              bfr                3004         1903         1894               2938        1904           1889
XI543              bfr                3197         1899         2919               2582        1900           457
XI544              bfr                2914         1893         323                3197        1890           1892
XI545              bfr                2997         1894         1888               2914        1889           1886
XI550              bfr                2745         1888         1887               2614        1886           1885
XI558              bfr                3140         1887         454                2637        1885           2818
XI560              bfr                2599         2550         1875               3205        1883           1884
XI561              bfr                3205         1882         1872               3130        1879           1881
XI571              bfr                2412         1878         1877               2906        456            1867
XI572              bfr                2889         398          1876               2412        399            1860
XI573              bfr                2906         1875         1856               2569        1884           1873
XI574              bfr                2569         1872         1859               3206        1881           1857
XI580              bfr                2702         1871         1870               2374        397            1845
XI581              bfr                3217         1877         1851               3112        1867           1868
XI582              bfr                2374         452          1865               2378        1864           1866
XI583              bfr                2378         1876         1844               3217        1860           1841
XI584              bfr                3076         1859         1840               2598        1857           1858
XI585              bfr                3112         1856         1854               3076        1873           1855
XI587              bfr                2538         1865         812                2727        1866           810
XI588              bfr                2579         1852         853                3057        450            849
XI589              bfr                2353         1851         1848               2786        1868           1849
XI590              bfr                3057         1870         1846               2538        1845           1847
XI591              bfr                2727         1844         793                2353        1841           1843
XI592              bfr                2362         1840         1838               2358        1858           1839
XI593              bfr                2786         1854         1836               2362        1855           1837
XI594              bfr                3111         1832         1833               2909        1825           1834
XI595              bfr                2336         1832         1831               3111        1975           1822
XI596              bfr                1835         1830         1821               2801        1644           1829
XI597              bfr                2801         1828         1827               2333        1826           1819
XI598              bfr                2333         1828         1818               2336        1825           1816
XI599              bfr                2972         1833         1823               2946        1834           1812
XI600              bfr                3164         1831         1811               2972        1822           1809
XI601              bfr                2958         1821         1808               3083        1829           1805
XI602              bfr                3083         1827         1804               2316        1819           1802
XI603              bfr                2316         1818         1817               3164        1816           1801
XI604              bfr                2524         1823         1813               2805        1812           1814
XI605              bfr                2304         1811         1796               2524        1809           1810
XI606              bfr                3067         1808         1807               2296        1805           1791
XI607              bfr                2296         1804         1803               2489        1802           1789
XI608              bfr                2489         1817         1788               2304        1801           1786
XI609              bfr                3165         1813         1797               2288        1814           1798
XI610              bfr                2684         1796         1794               3165        1810           1795
XI611              bfr                1820         1807         1781               3087        1791           1793
XI612              bfr                3087         1803         1778               2986        1789           1790
XI613              bfr                2986         1788         1776               2684        1786           1787
XI614              bfr                2835         1797         1784               2868        1798           1771
XI615              bfr                3061         1794         1782               2835        1795           1783
XI616              bfr                2971         1781         1770               2873        1793           1780
XI617              bfr                2873         1778         1768               2693        1790           1777
XI618              bfr                2693         1776         1774               3061        1787           1775
XI619              bfr                3098         1784         1772               2823        1771           1763
XI620              bfr                3097         1782         1762               3098        1783           1761
XI621              bfr                1806         1770         1757               2237        1780           1756
XI622              bfr                2237         1768         1767               2999        1777           1754
XI623              bfr                2999         1774         1760               3097        1775           1766
XI624              bfr                3215         1772         1764               3004        1763           1751
XI625              bfr                2712         1762         1750               3215        1761           1749
XI626              bfr                2822         1760         1759               2712        1766           1740
XI627              bfr                1800         1757         1748               2610        1756           1744
XI628              bfr                2610         1767         1755               2822        1754           1742
XI629              bfr                2893         1764         1752               2997        1751           1753
XI630              bfr                2210         1750         1739               2893        1749           1734
XI631              bfr                3079         1748         1746               3141        1744           1747
XI632              bfr                3141         1755         1727               2927        1742           1743
XI633              bfr                2927         1759         1741               2210        1740           1728
XI634              bfr                2602         1739         1735               2966        1734           1736
XI635              bfr                1785         1746         1732               2198        1747           1733
XI636              bfr                2711         1741         1730               2602        1728           1731
XI637              bfr                2198         1727         1718               2711        1743           1726
XI638              bfr                2966         1752         1725               2745        1753           1722
XI639              bfr                2177         1725         314                3140        1722           1723
XI640              bfr                2191         1730         1721               3170        1731           1708
XI641              bfr                1779         1732         1720               2782        1733           1710
XI642              bfr                2782         1718         1716               2191        1726           1717
XI643              bfr                3170         1735         1707               2177        1736           1705
XI644              bfr                2525         1716         1713               3055        1717           1714
XI645              bfr                3086         1720         1711               2525        1710           1712
XI646              bfr                3055         1721         1704               2166        1708           1702
XI647              bfr                2166         1707         1706               2586        1705           1699
XI649              bfr                2879         1711         1696               2528        1712           1693
XI650              bfr                2810         1704         306                2692        1702           305
XI651              bfr                2528         1713         1698               2810        1714           1701
XI652              bfr                2692         1706         445                3218        1699           1700
XI654              bfr                3201         1698         1689               2591        1701           1697
XI655              bfr                2864         1696         1694               3201        1693           1695
XI661              bfr                1758         1694         1690               2496        1695           1691
XI662              bfr                2496         1689         444                2548        1697           3065
XI674              bfr                1906         1688         871                2579        1685           1687
XI681              bfr                2708         1830         1683               1835        1826           1684
XI682              bfr                2486         1683         1682               2958        1684           1678
XI683              bfr                2677         1682         1677               3067        1678           1679
XI684              bfr                1686         1677         1676               1820        1679           1672
XI685              bfr                2792         1676         1674               2971        1672           1675
XI686              bfr                2900         1674         1671               1806        1675           1669
XI687              bfr                2736         1671         1670               1800        1669           1666
XI688              bfr                1709         1670         1667               3079        1666           1665
XI689              bfr                1715         1667         1664               1785        1665           1660
XI690              bfr                1719         1664         1662               1779        1660           1663
XI691              bfr                2698         1662         1659               3086        1663           1657
XI692              bfr                2636         1659         1656               2879        1657           1658
XI693              bfr                2859         1656         1654               2864        1658           1652
XI694              bfr                2916         1654         1653               1758        1652           1648
XI695              bfr                3090         1653         1650               1738        1648           1651
XI696              bfr                1655         1650         3448               1745        1651           595
XI697              bfr                1638         1647         1645               2708        1644           1646
XI698              bfr                1547         1643         1615               2859        1641           1611
XI699              bfr                2706         1639         1643               2636        1640           1641
XI700              bfr                3017         1636         1639               2698        1637           1640
XI701              bfr                2603         1633         1636               1719        1635           1637
XI702              bfr                2850         1634         1633               1715        1630           1635
XI703              bfr                1612         1632         1634               1709        1629           1630
XI704              bfr                2544         1626         1632               2736        1628           1629
XI705              bfr                2497         1627         1626               2900        1624           1628
XI706              bfr                2675         1622         1627               2792        1623           1624
XI707              bfr                2713         1617         1622               1686        1618           1623
XI708              bfr                1582         1621         1617               2677        1616           1618
XI709              bfr                1577         1645         1621               2486        1646           1616
XI710              bfr                2647         1615         1613               2916        1611           1614
XI711              bfr                1561         1610         372                1655        1608           1609
XI712              bfr                2885         1613         1610               3090        1614           1608
XI713              bfr                1541         1647         1605               1638        1528           1606
XI714              bfr                1450         1601         1604               1547        1602           1574
XI715              bfr                1473         1603         1601               2706        1599           1602
XI716              bfr                1535         1597         1603               3017        1598           1599
XI717              bfr                1529         1594         1597               2603        1595           1598
XI718              bfr                1523         1591         1594               2850        1593           1595
XI719              bfr                2866         1592         1591               1612        1590           1593
XI720              bfr                1512         1587         1592               2544        1588           1590
XI721              bfr                1506         1584         1587               2497        1585           1588
XI722              bfr                2638         1586         1584               2675        1583           1585
XI723              bfr                2485         1580         1586               2713        1581           1583
XI724              bfr                2580         1578         1580               1582        1579           1581
XI725              bfr                3101         1605         1578               1577        1606           1579
XI726              bfr                2728         1604         1575               2647        1574           1576
XI727              bfr                1460         1570         1573               1561        1571           2360
XI728              bfr                2977         1575         1570               2885        1576           1571
XI729              bfr                1443         1531         1540               1541        1487           1569
XI730              bfr                1351         1565         1538               1450        1566           1568
XI731              bfr                1376         1562         1565               1473        1563           1566
XI732              bfr                1438         1564         1562               1535        1559           1563
XI733              bfr                1431         1556         1564               1529        1558           1559
XI734              bfr                1423         1557         1556               1523        1555           1558
XI735              bfr                1418         1554         1557               2866        1552           1555
XI736              bfr                1413         1549         1554               1512        1551           1552
XI737              bfr                1406         1550         1549               1506        1548           1551
XI738              bfr                1401         1545         1550               2638        1546           1548
XI739              bfr                1395         1542         1545               2485        1544           1546
XI740              bfr                1389         1543         1542               2580        1539           1544
XI741              bfr                1383         1540         1543               3101        1569           1539
XI742              bfr                1356         1538         1536               2728        1568           1537
XI743              bfr                1363         1532         223                1460        1533           1534
XI744              bfr                1368         1536         1532               2977        1537           1533
XI745              bfr                1345         1531         1502               1443        1528           1530
XI746              bfr                1254         1527         1500               1351        1526           1496
XI747              bfr                1279         1525         1527               1376        1524           1526
XI748              bfr                1338         1521         1525               1438        1522           1524
XI749              bfr                1332         1519         1521               1431        1520           1522
XI750              bfr                3119         1516         1519               1423        1517           1520
XI751              bfr                1321         1514         1516               1418        1515           1517
XI752              bfr                1313         1511         1514               1413        1513           1515
XI753              bfr                1307         1509         1511               1406        1510           1513
XI754              bfr                1302         1507         1509               1401        1508           1510
XI755              bfr                1296         1503         1507               1395        1505           1508
XI756              bfr                1292         1504         1503               1389        1501           1505
XI757              bfr                1286         1502         1504               1383        1530           1501
XI758              bfr                1260         1500         1493               1356        1496           1497
XI759              bfr                1267         1495         2359               1363        1492           1494
XI760              bfr                1273         1493         1495               1368        1497           1492
XI761              bfr                1248         1490         1488               1345        1487           1489
XI762              bfr                1157         1486         1459               1254        1485           1457
XI763              bfr                1182         1484         1486               1279        1481           1485
XI764              bfr                1241         1482         1484               1338        1480           1481
XI765              bfr                1236         1476         1482               1332        1477           1480
XI766              bfr                1230         1478         1476               3119        1475           1477
XI767              bfr                2751         1471         1478               1321        1472           1475
XI768              bfr                1217         1474         1471               1313        1470           1472
XI769              bfr                1213         1468         1474               1307        1469           1470
XI770              bfr                1206         1465         1468               1302        1466           1469
XI771              bfr                1201         1462         1465               1296        1463           1466
XI772              bfr                1195         1464         1462               1292        1461           1463
XI773              bfr                1187         1488         1464               1286        1489           1461
XI774              bfr                1163         1459         1453               1260        1457           1458
XI775              bfr                1168         1456         185                1267        1452           1455
XI776              bfr                1174         1453         1456               1273        1458           1452
XI777              bfr                1150         1490         1451               1248        1371           1421
XI778              bfr                1064         1447         1420               1157        1448           1449
XI779              bfr                2840         1444         1447               1182        1445           1448
XI780              bfr                1145         1446         1444               1241        1442           1445
XI781              bfr                1140         1439         1446               1236        1441           1442
XI782              bfr                3212         1440         1439               1230        1436           1441
XI783              bfr                1128         1433         1440               2751        1434           1436
XI784              bfr                1122         1435         1433               1217        1432           1434
XI785              bfr                1116         1428         1435               1213        1429           1432
XI786              bfr                3176         1430         1428               1206        1427           1429
XI787              bfr                1103         1426         1430               1201        1425           1427
XI788              bfr                3223         1424         1426               1195        1422           1425
XI789              bfr                1094         1451         1424               1187        1421           1422
XI79               bfr                1824         2379         1815               514         329            332
XI790              bfr                1069         1420         1419               1163        1449           1415
XI791              bfr                3211         1417         2346               1168        1416           2344
XI792              bfr                1083         1419         1417               1174        1415           1416
XI793              bfr                1058         1414         1412               1150        1411           1382
XI794              bfr                964          1407         1381               1064        1409           1410
XI795              bfr                990          1408         1407               2840        1405           1409
XI796              bfr                1052         1404         1408               1145        1403           1405
XI797              bfr                1046         1399         1404               1140        1400           1403
XI798              bfr                1039         1402         1399               3212        1397           1400
XI799              bfr                1033         1398         1402               1128        1396           1397
XI80               bfr                505          334          1842               3418        345            332
XI800              bfr                1027         1392         1398               1122        1394           1396
XI801              bfr                1024         1393         1392               1116        1391           1394
XI802              bfr                1016         1387         1393               3176        1388           1391
XI803              bfr                1011         1390         1387               1103        1385           1388
XI804              bfr                1005         1386         1390               3223        1384           1385
XI805              bfr                998          1412         1386               1094        1382           1384
XI806              bfr                970          1381         1380               1069        1410           1373
XI807              bfr                974          1374         1378               3211        1377           1379
XI808              bfr                981          1380         1374               1083        1373           1377
XI809              bfr                957          1414         1372               1058        1371           1342
XI81               bfr                514          3441         1815               505         351            336
XI810              bfr                2783         1370         1341               964         1367           1369
XI811              bfr                893          1365         1370               990         1366           1367
XI812              bfr                954          1361         1365               1052        1362           1366
XI813              bfr                944          1364         1361               1046        1360           1362
XI814              bfr                2789         1357         1364               1039        1358           1360
XI815              bfr                935          1359         1357               1033        1355           1358
XI816              bfr                2949         1353         1359               1027        1354           1355
XI817              bfr                923          1349         1353               1024        1350           1354
XI818              bfr                918          1352         1349               1016        1348           1350
XI819              bfr                910          1346         1352               1011        1347           1348
XI82               bfr                3418         2419         1842               2243        2073           336
XI820              bfr                905          1343         1346               1005        1344           1347
XI821              bfr                899          1372         1343               998         1342           1344
XI822              bfr                873          1341         1339               970         1369           1340
XI823              bfr                880          1335         183                974         1336           1337
XI824              bfr                884          1339         1335               981         1340           1336
XI825              bfr                863          1334         1333               957         1411           1303
XI826              bfr                764          1327         1330               2783        1328           1331
XI827              bfr                795          1329         1327               893         1326           1328
XI828              bfr                858          1325         1329               954         1324           1326
XI829              bfr                850          1322         1325               944         1323           1324
XI830              bfr                844          1318         1322               2789        1319           1323
XI831              bfr                836          1320         1318               935         1317           1319
XI832              bfr                832          1316         1320               2949        1315           1317
XI833              bfr                827          1314         1316               923         1311           1315
XI834              bfr                820          1308         1314               918         1310           1311
XI835              bfr                814          1309         1308               910         1306           1310
XI836              bfr                806          1304         1309               905         1305           1306
XI837              bfr                3143         1333         1304               899         1303           1305
XI838              bfr                773          1330         1300               873         1331           1301
XI839              bfr                782          1299         1298               880         1297           181
XI84               bfr                3295         2380         2379               3370        341            329
XI840              bfr                790          1300         1299               884         1301           1297
XI841              bfr                755          1334         1268               863         1295           1265
XI842              bfr                636          1291         1264               764         1293           1294
XI843              bfr                2655         1289         1291               795         1290           1293
XI844              bfr                746          1287         1289               858         1288           1290
XI845              bfr                2623         1284         1287               850         1285           1288
XI846              bfr                3122         1281         1284               844         1283           1285
XI847              bfr                2817         1282         1281               836         1280           1283
XI848              bfr                3062         1276         1282               832         1277           1280
XI849              bfr                2828         1278         1276               827         1275           1277
XI850              bfr                3189         1274         1278               820         1271           1275
XI851              bfr                2549         1272         1274               814         1270           1271
XI852              bfr                681          1269         1272               806         1266           1270
XI853              bfr                2964         1268         1269               3143        1265           1266
XI854              bfr                2718         1264         1259               773         1294           1263
XI855              bfr                2856         1262         2306               782         1258           1261
XI856              bfr                2952         1259         1262               790         1263           1258
XI857              bfr                627          1218         1256               755         1177           1257
XI858              bfr                2503         1255         1226               636         1250           1224
XI859              bfr                2562         1251         1255               2655        1249           1250
XI86               bfr                547          2448         334                523         2449           345
XI860              bfr                618          1246         1251               746         1247           1249
XI861              bfr                611          1243         1246               2623        1244           1247
XI862              bfr                604          1245         1243               3122        1242           1244
XI863              bfr                2622         1239         1245               2817        1240           1242
XI864              bfr                586          1237         1239               3062        1238           1240
XI865              bfr                3116         1234         1237               2828        1235           1238
XI866              bfr                3033         1231         1234               3189        1232           1235
XI867              bfr                2514         1233         1231               2549        1229           1232
XI868              bfr                2541         1227         1233               681         1228           1229
XI869              bfr                3120         1256         1227               2964        1257           1228
XI870              bfr                2513         1226         1222               2718        1224           1219
XI871              bfr                3005         1220         1223               2856        1221           2286
XI872              bfr                2890         1222         1220               2952        1219           1221
XI873              bfr                3150         1218         1189               627         1295           1186
XI874              bfr                423          1216         1185               2503        1214           1215
XI875              bfr                440          1210         1216               2562        1211           1214
XI876              bfr                491          1212         1210               618         1209           1211
XI877              bfr                2858         1208         1212               611         1205           1209
XI878              bfr                2937         1207         1208               604         1204           1205
XI879              bfr                2661         1202         1207               2622        1203           1204
XI88               bfr                3370         2434         3441               547         421            351
XI880              bfr                3158         1198         1202               586         1199           1203
XI881              bfr                470          1200         1198               3116        1197           1199
XI882              bfr                465          1193         1200               3033        1196           1197
XI883              bfr                2996         1190         1193               2514        1192           1196
XI884              bfr                2512         1191         1190               2541        1188           1192
XI885              bfr                2564         1189         1191               3120        1186           1188
XI886              bfr                2491         1185         1184               2513        1215           1180
XI887              bfr                2519         1183         2278               3005        1181           2275
XI888              bfr                2590         1184         1183               2890        1180           1181
XI889              bfr                2609         1141         1178               3150        1177           1179
XI890              bfr                3115         1176         1148               423         1173           1175
XI891              bfr                3010         1172         1176               440         1170           1173
XI892              bfr                2710         1171         1172               491         1169           1170
XI893              bfr                406          1166         1171               2858        1167           1169
XI894              bfr                2539         1164         1166               2937        1165           1167
XI895              bfr                2793         1160         1164               2661        1162           1165
XI896              bfr                3225         1161         1160               3158        1159           1162
XI897              bfr                386          1155         1161               470         1156           1159
XI898              bfr                2871         1158         1155               465         1153           1156
XI899              bfr                3053         1154         1158               2996        1152           1153
XI90               bfr                523          3438         2419               2322        376            2073
XI900              bfr                3043         1151         1154               2512        1149           1152
XI901              bfr                3187         1178         1151               2564        1179           1149
XI902              bfr                2492         1148         1143               2491        1175           1147
XI903              bfr                2536         1146         1144               2519        1142           24
XI904              bfr                3190         1143         1146               2590        1147           1142
XI905              bfr                2816         1141         1113               2609        3499           1111
XI906              bfr                3041         1139         1110               3115        1138           1107
XI907              bfr                3175         1133         1139               3010        1137           1138
XI908              bfr                2739         1136         1133               2710        1132           1137
XI909              bfr                2483         1129         1136               406         1131           1132
XI91               bfr                2134         2421         2380               3356        3414           341
XI910              bfr                2594         1130         1129               2539        1127           1131
XI911              bfr                3160         1125         1130               2793        1126           1127
XI912              bfr                2668         1121         1125               3225        1124           1126
XI913              bfr                3002         1123         1121               386         1120           1124
XI914              bfr                2920         1119         1123               2871        1118           1120
XI915              bfr                2504         1117         1119               3053        1115           1118
XI916              bfr                3226         1114         1117               3043        1112           1115
XI917              bfr                2687         1113         1114               3187        1111           1112
XI918              bfr                2969         1110         1106               2492        1107           1108
XI919              bfr                226          1104         2240               2536        1105           2239
XI92               bfr                2161         3347         2421               3429        3369           3414
XI920              bfr                2807         1106         1104               3190        1108           1105
XI921              bfr                2910         1066         1101               2816        3496           1102
XI922              bfr                2717         1101         1100               2687        1102           1098
XI923              bfr                3114         1100         1099               3226        1098           1096
XI924              bfr                3121         1099         1097               2504        1096           1093
XI925              bfr                193          1097         1092               2920        1093           1095
XI926              bfr                186          1092         1091               3002        1095           1090
XI927              bfr                195          1091         1089               2668        1090           1085
XI928              bfr                194          1089         1086               3160        1085           1087
XI929              bfr                196          1086         1084               2594        1087           1082
XI93               bfr                3428         2441         3347               3337        453            3369
XI930              bfr                189          1084         1081               2483        1082           1079
XI931              bfr                188          1081         1078               2739        1079           1080
XI932              bfr                3139         1078         1076               3175        1080           1077
XI933              bfr                190          1076         1072               3041        1077           1073
XI934              bfr                2884         1072         1071               2969        1073           1068
XI935              bfr                3089         1071         1067               2807        1068           1070
XI936              bfr                192          1067         2258               226         1070           2257
XI937              bfr                3173         1066         1065               2910        3499           1036
XI938              bfr                200          1061         1063               190         1062           1032
XI939              bfr                197          1059         1061               3139        1060           1062
XI94               bfr                3444         2392         2441               235         3416           453
XI940              bfr                205          1056         1059               188         1057           1060
XI941              bfr                203          1053         1056               189         1055           1057
XI942              bfr                202          1054         1053               196         1051           1055
XI943              bfr                2956         1048         1054               194         1050           1051
XI944              bfr                2908         1049         1048               195         1047           1050
XI945              bfr                187          1043         1049               186         1045           1047
XI946              bfr                3015         1044         1043               193         1042           1045
XI947              bfr                227          1041         1044               3121        1040           1042
XI948              bfr                224          1037         1041               3114        1038           1040
XI949              bfr                2615         1065         1037               2717        1036           1038
XI95               bfr                3417         2385         2392               3446        3310           3416
XI950              bfr                229          1063         1034               2884        1032           1035
XI951              bfr                228          1031         1029               192         1028           1030
XI952              bfr                214          1034         1031               3089        1035           1028
XI953              bfr                201          987          1000               3173        3496           997
XI954              bfr                3034         1025         996                200         1026           993
XI955              bfr                3156         1022         1025               197         1023           1026
XI956              bfr                3224         1019         1022               205         1021           1023
XI957              bfr                204          1020         1019               203         1018           1021
XI958              bfr                2941         1017         1020               202         1014           1018
XI959              bfr                2877         1012         1017               2956        1013           1014
XI96               bfr                3440         2193         2385               3433        2430           3310
XI960              bfr                208          1009         1012               2908        1010           1013
XI961              bfr                211          1006         1009               187         1007           1010
XI962              bfr                242          1008         1006               3015        1004           1007
XI963              bfr                241          1001         1008               227         1003           1004
XI964              bfr                240          1002         1001               224         999            1003
XI965              bfr                244          1000         1002               2615        997            999
XI966              bfr                243          996          994                229         993            995
XI967              bfr                2762         988          991                228         989            992
XI968              bfr                2694         994          988                214         995            989
XI969              bfr                2924         987          985                201         3500           986
XI97               bfr                115          2233         2448               3335        2395           2449
XI970              bfr                212          984          982                3034        979            983
XI971              bfr                219          980          984                3156        978            979
XI972              bfr                218          977          980                3224        976            978
XI973              bfr                217          975          977                204         972            976
XI974              bfr                3193         973          975                2941        971            972
XI975              bfr                220          968          973                2877        969            971
XI976              bfr                3056         966          968                208         967            969
XI977              bfr                3066         962          966                211         963            967
XI978              bfr                246          965          962                242         961            963
XI979              bfr                250          960          965                241         959            961
XI98               bfr                301          2397         2233               273         2263           2395
XI980              bfr                248          958          960                240         956            959
XI981              bfr                3006         985          958                244         986            956
XI982              bfr                253          982          950                243         983            955
XI983              bfr                232          948          951                2762        949            952
XI984              bfr                231          950          948                2694        955            949
XI985              bfr                230          947          945                2924        3497           946
XI986              bfr                2618         941          919                212         942            915
XI987              bfr                3074         943          941                219         939            942
XI988              bfr                2896         940          943                218         938            939
XI989              bfr                237          936          940                217         937            938
XI99               bfr                3375         2425         2397               283         2386           2263
XI990              bfr                236          932          936                3193        934            937
XI991              bfr                239          933          932                220         931            934
XI992              bfr                2794         928          933                3056        929            931
XI993              bfr                238          930          928                3066        927            929
XI994              bfr                247          924          930                246         925            927
XI995              bfr                251          926          924                250         922            925
XI996              bfr                249          920          926                248         921            922
XI997              bfr                3199         945          920                3006        946            921
XI998              bfr                254          919          916                253         915            917
XI999              bfr                252          911          913                232         912            914
XI11               maj_bbb            2141         2500         2381               2388        2534           2164                   486   1919
XI12               maj_bbb            2370         2213         2221               1225        407            3493                   2367  479
XI153              maj_bbb            725          698          553                3448        635            767                    595   777
XI162              maj_bbb            701          651          638                409         2373           775                    408   2372
XI171              maj_bbb            621          564          538                3334        261            554                    477   2369
XI197              maj_bbb            697          739          362                476         741            668                    3330  1729
XI208              maj_bbb            364          691          509                3329        1681           347                    3328  1673
XI213              maj_bbb            308          709          206                3284        2349           702                    474   3327
XI22               maj_bbb            1968         2307         2022               485         2034           2348                   3346  1964
XI223              maj_bbb            737          641          142                3149        472            160                    3318  473
XI23               maj_bbb            2382         1737         1799               3342        482            3490                   2147  383
XI243              maj_bbb            67           57           615                686         1620           65                     140   624
XI33               maj_bbb            2194         2103         1375               3365        2273           3487                   487   2329
XI34               maj_bbb            2551         2314         2252               422         483            1619                   3279  2453
XI396              maj_bbb            3026         3322         3309               469         158            2540                   468   157
XI408              maj_bbb            2671         3315         3306               2720        467            3313                   495   2121
XI413              maj_bbb            3161         2632         3214               2144        2829           3305                   466   162
XI423              maj_bbb            3131         3289         2955               420         2113           3288                   419   2110
XI438              maj_bbb            2883         3270         2646               462         2083           2729                   418   2079
XI525              maj_bbb            2860         2641         2932               1942        116            2954                   461   2798
XI540              maj_bbb            2556         2757         2715               1910        120            2897                   2881  2803
XI547              maj_bbb            3011         2724         2730               459         1882           2691                   417   1879
XI555              maj_bbb            2776         2530         3184               2919        3191           2529                   457   2838
XI562              maj_bbb            2800         2533         2589               416         1878           2599                   415   456
XI568              maj_bbb            2870         2857         3132               454         135            2440                   2818  2703
XI575              maj_bbb            2581         2487         2732               414         452            2889                   451   1864
XI586              maj_bbb            2058         2645         1971               3096        1852           2702                   446   450
XI658              maj_bbb            3179         2065         2481               445         2970           2089                   1700  108
XI670              maj_bbb            2963         2733         2826               444         102            3144                   3065  103
XI677              maj_bbb            2842         2555         3185               2876        442            1906                   410   872
XI164              maj_bbi            600          518          542                722         284            638                    689   3269
XI18               maj_bbi            1978         2080         1997               2170        2458           2221                   1880  2457
XI206              maj_bbi            727          352          333                670         404            538                    713   566
XI216              maj_bbi            548          216          580                562         191            206                    607   525
XI225              maj_bbi            35           711          12                 723         3387           142                    1649  3382
XI29               maj_bbi            2118         2256         2201               1945        3349           1799                   2420  392
XI41               maj_bbi            2300         1560         1895               2339        3276           2252                   2650  2450
XI411              maj_bbi            3311         3307         3301               152         2921           3306                   153   403
XI427              maj_bbi            3171         3203         3080               172         2106           2955                   3093  2105
XI440              maj_bbi            2846         2891         2779               2785        2078           2646                   179   2076
XI552              maj_bbi            2488         2917         2584               131         2550           2730                   3125  1883
XI565              maj_bbi            2597         2895         2494               3027        398            2589                   137   399
XI578              maj_bbi            2957         2390         2384               146         1871           2732                   2628  397
XI668              maj_bbi            2571         2627         2482               100         1688           1971                   101   1685
XI678              maj_bbi            2775         1853         2833               3042        3147           3185                   105   395
XI14               maj_bib            2621         3373         2427               2663        2170           2213                   2605  1880
XI160              maj_bib            762          662          532                1869        722            651                    533   689
XI203              maj_bib            402          377          588                1765        670            564                    639   713
XI214              maj_bib            295          493          688                748         562            709                    1692  607
XI224              maj_bib            779          744          614                1661        723            641                    1668  1649
XI25               maj_bib            1680         2069         2325               2709        1945           1737                   2282  2420
XI36               maj_bib            2204         1498         1437               1863        2339           2314                   2447  2650
XI406              maj_bib            3319         3316         2750               151         152            3315                   3009  153
XI425              maj_bib            3293         3285         2902               2754        172            3289                   3084  3093
XI439              maj_bib            2848         2747         2629               2809        2785           3270                   2820  179
XI548              maj_bib            2983         2673         2626               2918        131            2724                   3025  3125
XI564              maj_bib            2748         3037         2624               126         3027           2533                   2831  137
XI576              maj_bib            2554         2625         3196               133         146            2487                   2961  2628
XI665              maj_bib            2802         2527         3020               112         100            2645                   2608  101
XI675              maj_bib            2516         2600         2619               2930        3042           2555                   114   105
XI13               maj_ibb            2431         1891         2518               572         2663           2370                   381   2605
XI155              maj_ibb            717          690          520                3447        1869           701                    292   533
XI199              maj_ibb            738          396          551                437         1765           621                    2925  639
XI209              maj_ibb            789          527          774                2787        748            308                    674   1692
XI219              maj_ibb            561          659          37                 2746        1661           737                    3297  1668
XI24               maj_ibb            2011         2042         1958               671         2709           2382                   384   2282
XI35               maj_ibb            2309         2508         2452               439         1863           2551                   438   2447
XI398              maj_ibb            3325         3168         3155               2774        151            2671                   435   3009
XI415              maj_ibb            3051         3292         2660               344         2754           3131                   342   3084
XI429              maj_ibb            3001         2553         2749               2701        2809           2883                   432   2820
XI541              maj_ibb            2773         2799         2657               431         2918           3011                   327   3025
XI556              maj_ibb            2758         2522         2547               321         126            2800                   429   2831
XI569              maj_ibb            2825         3102         3136               428         133            2581                   2752  2961
XI660              maj_ibb            3177         3077         2568               304         112            2058                   303   2608
XI672              maj_ibb            2654         2922         3172               426         2930           2842                   298   114
XI1                or_bb              2179         2229         2111               480         3494           645                    1075
XIsum0             sink               22           3392         3291               3271        0
XIsum1             sink               3383         3294         3392               3321        3271
XIsum10            sink               3044         2470         2467               2466        2468
XIsum11            sink               174          2472         2470               2469        2466
XIsum12            sink               176          2474         2472               2475        2469
XIsum13            sink               165          2476         2474               2473        2475
XIsum14            sink               159          2478         2476               2479        2473
XIsum15            sink               154          2480         2478               2477        2479
XIsum16            sink               257          0            2480               3105        2477
XIsum2             sink               31           3402         3294               3380        3321
XIsum3             sink               3340         3126         3402               3282        3380
XIsum4             sink               33           3353         3126               3355        3282
XIsum5             sink               3333         3409         3353               3384        3355
XIsum6             sink               3401         3283         3409               3331        3384
XIsum7             sink               3228         2464         3283               3406        3331
XIsum8             sink               3024         2465         2464               2463        3406
XIsum9             sink               184          2467         2465               2468        2463
XI10               spl2               2243         389          560                1930        388            3275                   2393
XI1199             spl2               2393         2276         560                2225        2283           645                    3445
XI1200             spl2               2460         2093         2276               2143        2031           2283                   1994
XI189              spl2               478          372          371                725         1609           3021                   706
XI19               spl2               3491         379          3134               2141        198            378                    2249
XI193              spl2               455          371          367                698         3021           366                    735
XI195              spl2               433          369          2973               697         209            684                    412
XI196              spl2               668          367          437                553         366            2925                   768
XI20               spl2               3492         3134         581                2500        378            2402                   2127
XI201              spl2               788          2973         365                739         684            361                    382
XI204              spl2               82           728          2882               364         156            2863                   320
XI207              spl2               347          365          2787               362         361            674                    338
XI21               spl2               2284         581          687                2381        2402           1135                   2054
XI211              spl2               71           2882         360                691         2863           359                    631
XI218              spl2               65           360          2746               509         359            3297                   753
XI242              spl2               3442         136          356                67          3213           2854                   732
XI245              spl2               3424         356          494                57          2854           673                    45
XI248              spl2               3487         494          439                615         673            438                    13
XI30               spl2               3488         2174         2343               1968        2429           3047                   1874
XI31               spl2               3489         2343         3230               2307        3047           1918                   2633
XI32               spl2               2164         3230         572                2022        1918           381                    2526
XI395              spl2               2953         2149         350                3026        2874           348                    3323
XI401              spl2               2950         350          343                3322        348            349                    3220
XI409              spl2               3127         346          340                3161        3142           337                    3148
XI412              spl2               3305         343          344                3309        349            342                    3304
XI416              spl2               3064         340          3088               2632        337            339                    3286
XI42               spl2               3485         393          3022               2194        88             374                    1912
XI428              spl2               2954         3088         2701               3214        339            432                    3278
XI43               spl2               3486         3022         3235               2103        374            528                    2377
XI44               spl2               2348         3235         671                1375        528            384                    2410
XI524              spl2               3103         1936         2821               2860        2679           335                    2944
XI532              spl2               2731         2821         328                2641        335            325                    2855
XI537              spl2               2813         331          324                2556        3180           330                    2995
XI539              spl2               2897         328          431                2932        325            327                    2790
XI546              spl2               2582         324          319                2757        330            318                    2699
XI551              spl2               2614         323          316                2776        1892           322                    2824
XI554              spl2               2529         319          321                2715        318            429                    2595
XI559              spl2               2637         316          317                2530        322            315                    2484
XI567              spl2               2440         317          428                3184        315            2752                   3071
XI648              spl2               2586         314          311                2870        1723           313                    2157
XI653              spl2               3218         311          312                2857        313            310                    2122
XI656              spl2               2591         306          309                3179        305            300                    3039
XI657              spl2               2089         312          304                3132        310            303                    2511
XI663              spl2               2548         309          302                2065        300            297                    2596
XI666              spl2               1738         1690         294                2963        1691           299                    3078
XI669              spl2               3144         302          426                2481        297            298                    2797
XI673              spl2               1745         294          296                2733        299            293                    3118
XI680              spl2               767          296          3447               2826        293            292                    1850
XI8                spl2               2322         2417         389                2640        2418           388                    2460
XI15               spl3L              2127         2266         2396               1891        2423           2558                   3373  2080
XI154              spl3L              706          635          1792               717         777            730                    762   600
XI16               spl3L              2249         2534         2266               2431        1919           2423                   2621  1978
XI161              spl3L              735          1792         705                690         730            2471                   662   518
XI163              spl3L              768          705          3334               520         2471           477                    532   542
XI17               spl3L              2054         2396         480                2518        2558           1075                   2427  1997
XI198              spl3L              412          741          663                738         1729           791                    402   727
XI202              spl3L              382          663          1769               396         791            1773                   377   352
XI205              spl3L              338          1769         3284               551         1773           474                    588   333
XI210              spl3L              320          1681         634                789         1673           1703                   295   548
XI215              spl3L              631          634          597                527         1703           1724                   493   216
XI217              spl3L              753          597          3149               774         1724           3318                   688   580
XI244              spl3L              732          1620         1625               561         624            1631                   779   35
XI246              spl3L              45           1625         582                659         1631           1642                   744   711
XI247              spl3L              13           582          422                37          1642           3279                   614   12
XI26               spl3L              2633         2261         1953               2042        2682           2563                   2069  2256
XI27               spl3L              1874         2034         2261               2011        1964           2682                   1680  2118
XI28               spl3L              2526         1953         1225               1958        2563           2367                   2325  2201
XI37               spl3L              2377         2456         2356               2508        2573           2416                   1498  1560
XI38               spl3L              1912         2273         2456               2309        2329           2573                   2204  2300
XI39               spl3L              2410         2356         3342               2452        2416           2147                   1437  1895
XI397              spl3L              3323         158          2898               3325        157            2934                   3319  3311
XI407              spl3L              3220         2898         2985               3168        2934           148                    3316  3307
XI410              spl3L              3304         2985         420                3155        148            419                    2750  3301
XI414              spl3L              3148         2829         3222               3051        162            163                    3293  3171
XI424              spl3L              3286         3222         3029               3292        163            169                    3285  3203
XI426              spl3L              3278         3029         462                2660        169            418                    2902  3080
XI526              spl3L              2944         116          117                3001        2798           2778                   2848  2846
XI533              spl3L              2855         117          125                2553        2778           123                    2747  2891
XI538              spl3L              2790         125          459                2749        123            417                    2629  2779
XI542              spl3L              2995         120          121                2773        2803           119                    2983  2488
XI549              spl3L              2699         121          3146               2799        119            128                    2673  2917
XI553              spl3L              2595         3146         416                2657        128            415                    2626  2584
XI557              spl3L              2824         3191         127                2758        2838           3181                   2748  2597
XI563              spl3L              2484         127          139                2522        3181           2915                   3037  2895
XI566              spl3L              3071         139          414                2547        2915           451                    2624  2494
XI570              spl3L              2157         135          134                2825        2703           3023                   2554  2957
XI577              spl3L              2122         134          144                3102        3023           143                    2625  2390
XI579              spl3L              2511         144          3096               3136        143            446                    3196  2384
XI659              spl3L              3039         2970         3219               3177        108            3007                   2802  2571
XI664              spl3L              2596         3219         98                 3077        3007           97                     2527  2627
XI667              spl3L              2797         98           2876               2568        97             410                    3020  2482
XI671              spl3L              3078         102          2744               2654        103            2832                   2516  2775
XI676              spl3L              3118         2744         104                2922        2832           2905                   2600  1853
XI679              spl3L              1850         104          409                3172        2905           408                    2619  2833
*end of top cell   16bit_RCA_ene_opt


.tran              {{t_step}}ps       {{end}}ps    {{begin}}ps  {{t_step}}ps
.FiLE              {{out_file_name}}
.print             i(Rac1)
*vac1_tot
.print             nodev              3497         0

.print             i(Rac2)
*vac2_tot
.print             nodev              3500         0

*vac1_DUT
.print             nodev              3496         3495
*vac2_DUT
.print             nodev              3499         3498