.model             jjmod                     jj(Rtype=1,  Vg=2.8mV,    Cap=0.064pF,  R0=100ohm,  Rn=17ohm,      Icrit=0.1mA)


.subckt            boost2_4_f4               1            2            3             54          55             56                     57    58    59
*inst name         cell_name                 a            din          dout          q1          q2             q3                     q4    xin   xout
B1                 15                        0            jjmod        area=0.5
B1a                51                        0            jjmod        area=0.5
B1b                19                        0            jjmod        area=0.5
B1c                22                        0            jjmod        area=0.5
B1d                30                        0            jjmod        area=0.5
B2                 34                        0            jjmod        area=0.5
B2a                18                        0            jjmod        area=0.5
B2b                9                         0            jjmod        area=0.5
B2c                20                        0            jjmod        area=0.5
B2d                28                        0            jjmod        area=0.5
Kd1                Ld                        L1           -0.133
Kd1a               Lda                       L1a          -0.133
Kd1b               Ldb                       L1b          -0.133
Kd1c               Ldc                       L1c          -0.133
Kd1d               Ldd                       L1d          -0.133
Kd2                Ld                        L2           -0.133
Kd2a               Lda                       L2a          -0.133
Kd2b               Ldb                       L2b          -0.133
Kd2c               Ldc                       L2c          -0.133
Kd2d               Ldd                       L2d          -0.133
Kdouta             Lda                       Louta        0.0
Kdoutb             Ldb                       Loutb        0.0
Kdoutc             Ldc                       Loutc        0.0
Kdoutd             Ldd                       Loutd        0.0
Kdqa               Lda                       Lqa          0.0
Kdqb               Ldb                       Lqb          0.0
Kdqc               Ldc                       Lqc          0.0
Kdqd               Ldd                       Lqd          0.0
Kouta              Lqa                       Louta        -0.495
Koutb              Lqb                       Loutb        -0.495
Koutd              Lqd                       Loutd        -0.495
Kqoutc             Lqc                       Loutc        -0.495
Kx1                Lx                        L1           -0.186
Kx1a               Lxa                       L1a          -0.186
Kx1b               Lxb                       L1b          -0.186
Kx1c               Lxc                       L1c          -0.186
Kx1d               Lxd                       L1d          -0.186
Kx2                Lx                        L2           -0.186
Kx2a               Lxa                       L2a          -0.186
Kx2b               Lxb                       L2b          -0.186
Kx2c               Lxc                       L2c          -0.186
Kx2d               Lxd                       L2d          -0.186
Kxd                Lx                        Ld           0.19
Kxda               Lxa                       Lda          0.19
Kxdb               Lxb                       Ldb          0.19
Kxdc               Lxc                       Ldc          0.19
Kxdd               Lxd                       Ldd          0.19
Kxouta             Lxa                       Louta        0.0
Kxoutb             Lxb                       Loutb        0.0
Kxoutc             Lxc                       Loutc        0.0
Kxoutd             Lxd                       Loutd        0.0
Kxqa               Lxa                       Lqa          0.0
Kxqb               Lxb                       Lqb          0.0
Kxqc               Lxc                       Lqc          0.0
Kxqd               Lxd                       Lqd          0.0
L1                 45                        15           1.59pH
L1a                50                        51           1.59pH
L1b                49                        19           1.59pH
L1c                40                        22           1.59pH
L1d                48                        30           1.59pH
L2                 34                        45           1.59pH
L2a                18                        50           1.59pH
L2b                9                         49           1.59pH
L2c                20                        40           1.59pH
L2d                28                        48           1.59pH
Ld                 2                         6            7.45pH
Lda                6                         5            7.45pH
Ldb                5                         41           7.45pH
Ldc                41                        46           7.45pH
Ldd                46                        3            7.45pH
Lin                1                         45           1.23pH
Lina               4                         50           3.4pH
Linb               4                         49           3.0pH
Linc               4                         40           3.0pH
Lind               4                         48           3.4pH
Louta              25                        54           31.2pH
Loutb              17                        55           31.2pH
Loutc              38                        56           31.2pH
Loutd              47                        57           31.2pH
Lq                 45                        4            9.96pH
Lqa                50                        53           7.92pH
Lqb                49                        24           7.92pH
Lqc                40                        26           7.92pH
Lqd                48                        32           7.92pH
Lx                 58                        7            7.4pH
Lxa                7                         8            7.4pH
Lxb                8                         16           7.4pH
Lxc                16                        43           7.4pH
Lxd                43                        59           7.4pH
R1a                25                        0            1e-12ohm
R1b                17                        0            1e-12ohm
R4                 53                        0            1e-12ohm
R5                 24                        0            1e-12ohm
R6                 38                        0            1e-12ohm
R7                 26                        0            1e-12ohm
R8                 47                        0            1e-12ohm
R9                 32                        0            1e-12ohm
.ends


.subckt            boost2_3_f3               1            2            3             41          42             43                     44    45
*inst name         cell_name                 a            din          dout          q1          q2             q3                     xin   xout
B1                 11                        0            jjmod        area=0.5
B1a                36                        0            jjmod        area=0.5
B1b                14                        0            jjmod        area=0.5
B1c                17                        0            jjmod        area=0.5
B2                 24                        0            jjmod        area=0.5
B2a                13                        0            jjmod        area=0.5
B2b                5                         0            jjmod        area=0.5
B2c                15                        0            jjmod        area=0.5
Kd1                Ld                        L1           -0.0644
Kd1a               Ld                        L1a          -0.0639
Kd1b               Ld                        L1b          -0.0662
Kd1c               Ld                        L1c          -0.066
Kd2                Ld                        L2           -0.0646
Kd2a               Ld                        L2a          -0.0653
Kd2b               Ld                        L2b          -0.0666
Kd2c               Ld                        L2c          -0.0642
Kdouta             Ld                        Louta        0.0007254
Kdoutb             Ld                        Loutb        0.0004117
Kdoutc             Ld                        Loutc        -0.001253
Kdq                Ld                        Lq           0.0
Kdqa               Ld                        Lqa          -0.0006276
Kdqb               Ld                        Lqb          -0.0005469
Kdqc               Ld                        Lqc          0.001507
Kdql               Ld                        Lql          0.0
Kdqr               Ld                        Lqr          0.0
Kouta              Lqa                       Louta        -0.493
Koutb              Lqb                       Loutb        -0.493
Koutc              Lqc                       Loutc        -0.493
Kx1                Lx                        L1           -0.0881
Kx1a               Lx                        L1a          -0.0893
Kx1b               Lx                        L1b          -0.0909
Kx1c               Lx                        L1c          -0.0907
Kx2                Lx                        L2           -0.0885
Kx2a               Lx                        L2a          -0.0903
Kx2b               Lx                        L2b          -0.0908
Kx2c               Lx                        L2c          -0.0894
Kxd                Lx                        Ld           0.177
Kxouta             Lx                        Louta        0.0003079
Kxoutb             Lx                        Loutb        -9.704e-05
Kxoutc             Lx                        Loutc        -0.0003689
Kxq                Lx                        Lq           0.0
Kxqa               Lx                        Lqa          -0.0003187
Kxqb               Lx                        Lqb          -0.0003226
Kxqc               Lx                        Lqc          0.0008805
Kxql               Lx                        Lql          0.0
Kxqr               Lx                        Lqr          0.0
L1                 31                        11           1.58pH
L1a                34                        36           1.49pH
L1b                32                        14           1.49pH
L1c                29                        17           1.49pH
L2                 24                        31           1.58pH
L2a                13                        34           1.49pH
L2b                5                         32           1.49pH
L2c                15                        29           1.49pH
Ld                 2                         3            36.97pH
Lin                1                         31           2.03pH
Lina               33                        34           1.23pH
Linb               4                         32           1.37pH
Linc               37                        29           1.36pH
Louta              20                        41           31.1pH
Loutb              12                        42           31.1pH
Loutc              27                        43           31.1pH
Lq                 31                        35           7.76pH
Lqa                34                        39           7.9pH
Lqb                32                        19           7.89pH
Lqc                29                        21           7.91pH
Lql                35                        33           5.27pH
Lqr                40                        35           5.06pH
Lqrb               40                        4            0.19pH
Lqrc               40                        37           1.36pH
Lx                 44                        45           36.64pH
R1a                20                        0            1e-12ohm
R1b                12                        0            1e-12ohm
R4                 39                        0            1e-12ohm
R5                 19                        0            1e-12ohm
R6                 27                        0            1e-12ohm
R7                 21                        0            1e-12ohm
.ends


.subckt            branch3                   1            2            3             4
*inst name         cell_name                 a            b            c             d
Lip                7                         4            0.312pH
Lp1                1                         6            11.8pH
Lp2                2                         7            10.2pH
Lp3                3                         5            11.8pH
R0                 6                         7            1e-12ohm
R1                 5                         7            1e-12ohm
.ends


.subckt            bfr                       1            2            3             12          13             14
*inst name         cell_name                 a            din          dout          q           xin            xout
B1                 9                         0            jjmod        area=0.5
B2                 5                         0            jjmod        area=0.5
Kd1                Ld                        L1           -0.133
Kd2                Ld                        L2           -0.133
Kdout              Ld                        Lout         0.0
Kdq                Ld                        Lq           0.0
Kout               Lq                        Lout         -0.495
Kx1                Lx                        L1           -0.186
Kx2                Lx                        L2           -0.186
Kxd                Lx                        Ld           0.19
Kxout              Lx                        Lout         0.0
Kxq                Lx                        Lq           0.0
L1                 8                         9            1.59pH
L2                 5                         8            1.59pH
Ld                 2                         3            7.45pH
Lin                1                         8            1.23pH
Lout               6                         12           31.2pH
Lq                 8                         0            7.92pH
Lx                 13                        14           7.4pH
R1                 6                         0            1e-12ohm
.ends


.subckt            inv                       1            2            3             12          13             14
*inst name         cell_name                 a            din          dout          q           xin            xout
B1                 9                         0            jjmod        area=0.6
B2                 5                         0            jjmod        area=0.6
Kd1                Ld                        L1           -0.133
Kd2                Ld                        L2           -0.133
Kdout              Ld                        Lout         0.0
Kdq                Ld                        Lq           0.0
Kout               Lq                        Lout         0.432
Kx1                Lx                        L1           -0.186
Kx2                Lx                        L2           -0.186
Kxd                Lx                        Ld           0.19
Kxout              Lx                        Lout         0.0
Kxq                Lx                        Lq           0.0
L1                 8                         9            1.59pH
L2                 5                         8            1.59pH
Ld                 2                         3            7.44pH
Lin                1                         8            1.24pH
Lout               6                         12           31.0pH
Lq                 8                         0            6.49pH
Lx                 13                        14           7.39pH
R1                 6                         0            1e-12ohm
.ends


.subckt            maj_bbi                   1            2            3             4           5              13                     14    15
*inst name         cell_name                 a            b            c             din         dout           q                      xin   xout
XI0                bfr                       1            4            9             11          14             6
XI1                bfr                       2            9            12            7           6              8
XI3                branch3                   11           7            10            13
XI2                inv                       3            12           5             10          8              15
.ends


.subckt            const0                    1            2            11            12          13
*inst name         cell_name                 din          dout         q             xin         xout
B1                 8                         0            jjmod        area=0.5
B2                 4                         0            jjmod        area=0.5
Kd1                Ld                        L1           -0.128
Kd2                Ld                        L2           -0.135
Kdout              Ld                        Lout         -0.000253
Kdq                Ld                        Lq           -0.00468
Kout               Lq                        Lout         -0.495
Kx1                Lx                        L1           -0.185
Kx2                Lx                        L2           -0.189
Kxd                Lx                        Ld           0.193
Kxout              Lx                        Lout         -7.94e-05
Kxq                Lx                        Lq           -0.00421
L1                 7                         8            1.56pH
L2                 4                         7            1.66pH
Ld                 1                         2            7.49pH
Lout               5                         11           31.2pH
Lq                 7                         0            7.82pH
Lx                 12                        13           7.47pH
R1                 5                         0            1e-12ohm
.ends


.subckt            and_bb                    1            2            3             4           12             13                     14
*inst name         cell_name                 a            b            din           dout        q              xin                    xout
XI0                bfr                       1            3            8             9           13             5
XI2                bfr                       2            11           4             10          7              14
XI3                branch3                   9            6            10            12
XI1                const0                    8            11           6             5           7
.ends


.subckt            maj_bib                   1            2            3             4           5              13                     14    15
*inst name         cell_name                 a            b            c             din         dout           q                      xin   xout
XI0                bfr                       1            4            9             11          14             6
XI2                bfr                       3            7            5             10          8              15
XI3                branch3                   11           12           10            13
XI1                inv                       2            9            7             12          6              8
.ends


.subckt            maj_ibb                   1            2            3             4           5              13                     14    15
*inst name         cell_name                 a            b            c             din         dout           q                      xin   xout
XI1                bfr                       2            8            10            12          6              7
XI2                bfr                       3            10           5             9           7              15
XI3                branch3                   11           12           9             13
XI0                inv                       1            4            8             11          14             6
.ends


.subckt            maj_bbb                   1            2            3             4           5              13                     14    15
*inst name         cell_name                 a            b            c             din         dout           q                      xin   xout
XI0                bfr                       1            4            8             11          14             6
XI1                bfr                       2            8            10            12          6              7
XI2                bfr                       3            10           5             9           7              15
XI3                branch3                   11           12           9             13
.ends


.subckt            sink                      1            2            3             10          11
*inst name         cell_name                 a            din          dout          xin         xout
B1                 8                         0            jjmod        area=0.5
B2                 5                         0            jjmod        area=0.5
Kd1                Ld                        L1           -0.133
Kd2                Ld                        L2           -0.133
Kdq                Ld                        Lq           0.0
Kx1                Lx                        L1           -0.186
Kx2                Lx                        L2           -0.186
Kxd                Lx                        Ld           0.19
Kxq                Lx                        Lq           0.0
L1                 7                         8            1.59pH
L2                 5                         7            1.59pH
Ld                 2                         3            7.45pH
Lin                1                         7            1.23pH
Lq                 7                         0            7.92pH
Lx                 10                        11           7.4pH
.ends


.subckt            and_bi                    1            2            3             4           12             13                     14
*inst name         cell_name                 a            b            din           dout        q              xin                    xout
XI0                bfr                       1            3            8             9           13             5
XI3                branch3                   9            7            10            12
XI1                const0                    8            11           7             5           6
XI2                inv                       2            11           4             10          6              14
.ends


.subckt            and_ib                    1            2            3             4           12             13                     14
*inst name         cell_name                 a            b            din           dout        q              xin                    xout
XI2                bfr                       2            11           4             10          6              14
XI3                branch3                   9            8            10            12
XI1                const0                    7            11           8             5           6
XI0                inv                       1            3            7             9           13             5
.ends


.subckt            const1                    1            2            7             8           9
*inst name         cell_name                 din          dout         q             xin         xout
L1                 8                         4            0.01pH
L2                 6                         9            0.01pH
L3                 1                         3            0.01pH
L4                 5                         2            0.01pH
XI0                const0                    5            3            7             6           4
.ends


.subckt            or_bb                     1            2            3             4           12             13                     14
*inst name         cell_name                 a            b            din           dout        q              xin                    xout
XI0                bfr                       1            3            8             9           13             5
XI2                bfr                       2            11           4             10          6              14
XI3                branch3                   9            7            10            12
XI1                const1                    8            11           7             5           6
.ends


*this is top cell  8bit_RCA_ene_opt_booster
R0                 490                       795          1000.0ohm
R1                 618                       807          1000.0ohm
R10                785                       1036         1000.0ohm
R11                889                       1017         1000.0ohm
R12                878                       766          1000.0ohm
R13                872                       761          1000.0ohm
R14                876                       919          1000.0ohm
R15                902                       1011         1000.0ohm
R2                 526                       779          1000.0ohm
R3                 616                       447          1000.0ohm
R4                 762                       824          1000.0ohm
R5                 764                       811          1000.0ohm
R6                 595                       842          1000.0ohm
R7                 739                       698          1000.0ohm
R8                 897                       1027         1000.0ohm
R9                 778                       1002         1000.0ohm
Rac1               885                       1105         100000.0ohm
Rac2               866                       1108         100000.0ohm
Rdc1               905                       617          100000.0ohm
V29                902                       0            PWL          (0ps          0mv         20ps           {{input[0]}})
V30                872                       0            PWL          (0ps          0mv         20ps           {{input[1]}})
V31                889                       0            PWL          (0ps          0mv         20ps           {{input[2]}})
V32                778                       0            PWL          (0ps          0mv         20ps           {{input[3]}})
V33                739                       0            PWL          (0ps          0mv         20ps           {{input[4]}})
V34                764                       0            PWL          (0ps          0mv         20ps           {{input[5]}})
V35                616                       0            PWL          (0ps          0mv         20ps           {{input[6]}})
V36                618                       0            PWL          (0ps          0mv         20ps           {{input[7]}})
V37                490                       0            PWL          (0ps          0mv         20ps           {{input[8]}})
V38                526                       0            PWL          (0ps          0mv         20ps           {{input[9]}})
V39                762                       0            PWL          (0ps          0mv         20ps           {{input[10]}})
V40                595                       0            PWL          (0ps          0mv         20ps           {{input[11]}})
V41                897                       0            PWL          (0ps          0mv         20ps           {{input[12]}})
V42                785                       0            PWL          (0ps          0mv         20ps           {{input[13]}})
V43                878                       0            PWL          (0ps          0mv         20ps           {{input[14]}})
V44                876                       0            PWL          (0ps          0mv         20ps           {{input[15]}})
VDC                905                       0            PWL          (0ps          0mV         20ps           113000mV)
VAC1               885                       0            SIN          (0            81000mV     {{freq}}MEGHz  {{40+period|int/4}}ps  0)
VAC2               866                       0            SIN          (0            81000mV     {{freq}}MEGHz  40ps                   0)
XI333              and_bb                    529          468          737           441         771            506                    238
XI336              and_bi                    567          539          436           737         334            1057                   506
XI338              and_ib                    538          524          255           436         495            250                    1057
XI100              bfr                       956          995          748           1026        295            746
XI101              bfr                       126          931          995           483         226            295
XI102              bfr                       1009         972          931           1014        848            226
XI103              bfr                       965          283          808           147         835            805
XI104              bfr                       1018         827          283           247         922            835
XI105              bfr                       949          225          827           975         285            922
XI106              bfr                       217          800          225           956         982            285
XI107              bfr                       1038         271          800           126         273            982
XI108              bfr                       1019         594          271           1009        558            273
XI109              bfr                       943          979          242           84          241            757
XI110              bfr                       232          220          979           113         592            241
XI111              bfr                       237          1006         220           664         986            592
XI112              bfr                       1026         816          1006          34          817            986
XI113              bfr                       483          297          816           157         933            817
XI114              bfr                       1014         291          297           221         845            933
XI117              bfr                       1098         293          246           671         292            759
XI118              bfr                       671          849          249           843         289            774
XI119              bfr                       923          246          259           855         759            966
XI120              bfr                       743          243          854           923         248            852
XI121              bfr                       855          249          1041          930         774            987
XI122              bfr                       1101         960          667           743         1025           846
XI123              bfr                       1044         259          258           980         966            263
XI124              bfr                       980          1041         90            1004        987            257
XI125              bfr                       163          667          262           60          846            263
XI126              bfr                       1102         298          871           112         1045           250
XI127              bfr                       60           854          258           1044        852            282
XI128              bfr                       112          11           262           163         602            282
XI129              bfr                       34           793          65            279         791            264
XI130              bfr                       664          65           864           314         264            254
XI131              bfr                       84           268          666           215         267            78
XI132              bfr                       113          864          268           252         254            267
XI133              bfr                       555          773          287           624         240            227
XI134              bfr                       157          837          793           555         284            791
XI135              bfr                       314          184          918           424         286            260
XI136              bfr                       424          261          734           498         269            507
XI137              bfr                       221          45           837           521         46             284
XI138              bfr                       252          918          239           1099        260            229
XI139              bfr                       215          239          441           1100        229            238
XI140              bfr                       498          233          914           1097        913            419
XI141              bfr                       475          1040         233           1096        251            913
XI142              bfr                       672          566          904           1094        395            763
XI143              bfr                       680          904          663           1095        763            670
XI144              bfr                       668          236          277           672         228            580
XI145              bfr                       669          277          1032          680         580            809
XI146              bfr                       643          54           769           668         55             245
XI147              bfr                       596          275          266           643         348            296
XI148              bfr                       624          266          281           662         296            231
XI149              bfr                       662          769          1040          669         245            251
XI150              bfr                       372          281          261           475         231            269
XI151              bfr                       521          256          773           596         486            240
XI152              bfr                       279          287          184           372         227            286
XI373              bfr                       317          210          207           209         611            208
XI374              bfr                       205          740          193           204         203            581
XI375              bfr                       204          749          191           201         202            187
XI376              bfr                       199          365          196           198         200            197
XI377              bfr                       198          195          178           194         470            174
XI378              bfr                       194          193          173           190         581            192
XI379              bfr                       190          191          188           189         187            181
XI386              bfr                       185          186          482           183         430            478
XI387              bfr                       183          516          156           180         606            182
XI388              bfr                       180          196          179           177         197            543
XI389              bfr                       177          178          175           172         174            176
XI390              bfr                       172          173          166           171         192            170
XI391              bfr                       171          188          167           169         181            168
XI396              bfr                       165          428          142           162         742            140
XI397              bfr                       162          519          159           161         415            160
XI398              bfr                       161          482          520           155         478            158
XI399              bfr                       155          156          153           154         182            132
XI400              bfr                       154          179          131           152         543            151
XI401              bfr                       152          175          148           150         176            149
XI402              bfr                       150          166          146           145         170            487
XI403              bfr                       145          167          122           144         168            119
XI406              bfr                       843          142          513           139         140            141
XI407              bfr                       139          159          607           138         160            143
XI408              bfr                       138          520          135           134         158            136
XI409              bfr                       134          153          133           130         132            105
XI410              bfr                       130          131          127           129         151            128
XI411              bfr                       129          148          103           125         149            99
XI412              bfr                       125          146          98            121         487            570
XI413              bfr                       121          122          96            120         119            91
XI416              bfr                       930          513          116           118         141            541
XI417              bfr                       118          607          588           111         143            115
XI418              bfr                       111          135          86            109         136            110
XI419              bfr                       109          133          107           108         105            80
XI420              bfr                       108          127          123           104         128            542
XI421              bfr                       104          103          100           97          99             101
XI422              bfr                       97           98           74            94          570            501
XI423              bfr                       94           96           92            93          91             69
XI426              bfr                       1004         116          90            88          541            562
XI427              bfr                       88           588          83            87          115            257
XI428              bfr                       87           86           83            85          110            562
XI429              bfr                       85           107          534           79          80             81
XI430              bfr                       79           123          534           76          542            484
XI431              bfr                       76           100          72            75          101            81
XI432              bfr                       75           74           72            73          501            484
XI433              bfr                       73           92           70            71          69             1103
XI436              bfr                       68           472          66            474         114            67
XI437              bfr                       62           467          370           68          41             64
XI438              bfr                       63           37           566           62          38             395
XI439              bfr                       56           33           236           63          57             228
XI440              bfr                       50           28           54            56          29             55
XI441              bfr                       51           52           275           50          48             348
XI442              bfr                       47           22           256           51          586            486
XI443              bfr                       389          20           45            47          44             46
XI446              bfr                       42           43           472           1           10             114
XI447              bfr                       39           5            467           42          6              41
XI448              bfr                       35           40           37            39          36             38
XI449              bfr                       30           1088         33            35          1089           57
XI450              bfr                       31           1085         28            30          27             29
XI451              bfr                       23           577          52            31          82             48
XI452              bfr                       24           25           22            23          604            586
XI453              bfr                       21           1079         20            24          19             44
XI456              bfr                       17           18           15            792         1077           16
XI457              bfr                       12           77           731           17          1075           730
XI458              bfr                       13           53           43            12          8              10
XI459              bfr                       7            49           5             13          4              6
XI460              bfr                       1093         1068         40            7           1091           36
XI461              bfr                       1090         1065         1088          1093        564            1089
XI462              bfr                       1087         1061         1085          1090        1084           27
XI463              bfr                       1083         1056         577           1087        1058           82
XI464              bfr                       1082         1051         25            1083        1052           604
XI465              bfr                       416          1081         1079          1082        61             19
XI466              bfr                       1078         59           18            390         58             1077
XI467              bfr                       1071         380          77            1078        1074           1075
XI468              bfr                       1072         1073         53            1071        1030           8
XI469              bfr                       1070         26           49            1072        1069           4
XI470              bfr                       1066         545          1068          1070        1022           1091
XI471              bfr                       1062         1067         1065          1066        1064           564
XI472              bfr                       1059         1063         1061          1062        302            1084
XI473              bfr                       1053         1060         1056          1059        338            1058
XI474              bfr                       1054         1055         1051          1053        857            1052
XI475              bfr                       833          1050         1081          1054        1049           61
XI476              bfr                       431          427          851           316         455            753
XI477              bfr                       357          508          812           431         406            433
XI478              bfr                       1039         557          59            357         32             58
XI479              bfr                       452          454          380           1039        1034           1074
XI480              bfr                       422          510          1073          452         1028           1030
XI481              bfr                       461          990          26            422         400            1069
XI482              bfr                       347          398          545           461         1021           1022
XI483              bfr                       367          306          1067          347         515            1064
XI484              bfr                       1013         1086         1063          367         509            302
XI485              bfr                       460          1015         1060          1013        974            338
XI486              bfr                       459          369          427           336         14             455
XI487              bfr                       448          354          508           459         568            406
XI488              bfr                       998          404          557           448         9              32
XI489              bfr                       403          1076         454           998         957            1034
XI490              bfr                       992          480          510           403         3              1028
XI491              bfr                       993          339          990           992         1092           400
XI492              bfr                       335          556          398           993         358            1021
XI493              bfr                       300          305          306           335         981            515
XI494              bfr                       331          870          1086          300         351            509
XI495              bfr                       862          977          1015          331         457            974
XI496              bfr                       968          471          464           363         304            745
XI497              bfr                       969          554          597           968         936            725
XI498              bfr                       346          432          369           969         1080           14
XI499              bfr                       961          928          354           346         355            568
XI500              bfr                       962          376          404           961         377            9
XI501              bfr                       955          412          1076          962         569            957
XI502              bfr                       952          915          480           955         954            3
XI503              bfr                       953          912          339           952         453            1092
XI504              bfr                       399          906          556           953         907            358
XI505              bfr                       439          312          305           399         322            981
XI506              bfr                       941          942          471           2           940            304
XI507              bfr                       938          572          554           941         410            936
XI508              bfr                       929          572          432           938         940            1080
XI509              bfr                       401          456          928           929         410            355
XI510              bfr                       920          456          376           401         366            377
XI511              bfr                       921          522          412           920         579            569
XI512              bfr                       414          522          915           921         366            954
XI513              bfr                       908          413          912           414         579            453
XI514              bfr                       910          413          906           908         315            907
XI515              bfr                       886          349          312           910         473            322
XI516              bfr                       324          788          518           402         1104           1042
XI517              bfr                       402          392          880           411         1107           344
XI518              bfr                       411          392          890           888         473            891
XI519              bfr                       888          349          1024          886         315            397
XI520              bfr                       333          518          326           884         1042           883
XI521              bfr                       884          880          445           879         344            552
XI522              bfr                       879          890          977           874         891            457
XI523              bfr                       874          1024         870           439         397            351
XI524              bfr                       868          326          865           863         883            320
XI525              bfr                       863          445          860           862         552            383
XI526              bfr                       859          865          1050          311         320            1049
XI527              bfr                       311          860          1055          460         383            857
XI528              bfr                       698          612          429           697         841            278
XI529              bfr                       697          838          594           699         385            558
XI530              bfr                       699          997          972           700         847            848
XI531              bfr                       700          834          291           389         373            845
XI532              bfr                       842          309          612           711         303            841
XI533              bfr                       711          814          838           712         435            385
XI534              bfr                       712          359          997           709         996            847
XI535              bfr                       709          462          834           21          821            373
XI536              bfr                       701          775          831           833         830            820
XI537              bfr                       706          772          818           701         549            829
XI538              bfr                       705          589          815           706         442            813
XI539              bfr                       824          825          823           705         768            973
XI540              bfr                       707          831          462           416         820            821
XI541              bfr                       708          818          359           707         829            996
XI542              bfr                       710          815          814           708         813            435
XI543              bfr                       811          823          309           710         973            303
XI544              bfr                       807          458          437           723         384            806
XI545              bfr                       723          804          503           722         802            780
XI546              bfr                       722          789          368           704         801            783
XI547              bfr                       704          409          798           333         796            799
XI548              bfr                       795          617          458           703         1105           384
XI549              bfr                       703          794          804           715         1108           802
XI550              bfr                       715          794          789           714         1104           801
XI551              bfr                       714          788          409           324         1107           796
XI552              bfr                       716          798          777           868         799            786
XI553              bfr                       717          368          421           716         783            784
XI554              bfr                       719          503          469           717         780            782
XI555              bfr                       779          437          770           719         806            767
XI556              bfr                       718          777          775           859         786            830
XI557              bfr                       721          421          772           718         784            549
XI558              bfr                       720          469          589           721         782            442
XI559              bfr                       447          770          825           720         767            768
XI560              bfr                       209          533          608           505         1106           638
XI561              bfr                       505          533          644           535         328            634
XI562              bfr                       535          590          654           544         0              502
XI564              bfr                       747          608          651           593         638            574
XI566              bfr                       537          654          493           332         502            650
XI567              bfr                       593          644          630           537         634            583
XI568              bfr                       530          630          418           653         583            573
XI569              bfr                       653          493          517           645         650            477
XI570              bfr                       201          651          622           530         574            658
XI572              bfr                       628          418          599           499         573            494
XI573              bfr                       499          517          615           641         477            591
XI574              bfr                       189          622          640           628         658            476
XI576              bfr                       582          599          656           648         494            896
XI577              bfr                       648          615          633           639         591            479
XI578              bfr                       169          640          892           582         476            563
XI580              bfr                       625          656          585           525         896            511
XI581              bfr                       525          633          620           598         479            561
XI582              bfr                       144          892          489           625         563            626
XI584              bfr                       488          585          584           635         511            514
XI585              bfr                       635          620          877           621         561            875
XI586              bfr                       120          489          504           488         626            565
XI588              bfr                       637          584          613           657         514            642
XI589              bfr                       657          877          623           531         875            492
XI590              bfr                       93           504          497           637         565            614
XI593              bfr                       71           497          70            481         614            234
XI594              bfr                       649          623          587           632         492            234
XI595              bfr                       481          613          587           649         642            1103
XI83               bfr                       1011         211          1029          994         932            212
XI84               bfr                       919          946          211           971         216            932
XI85               bfr                       983          213          988           947         732            212
XI86               bfr                       440          218          213           425         214            732
XI87               bfr                       994          270          1029          983         219            758
XI88               bfr                       971          808          270           440         805            219
XI89               bfr                       947          265          988           822         1016           758
XI90               bfr                       425          242          265           790         757            1016
XI91               bfr                       761          222          946           965         999            216
XI92               bfr                       766          958          222           1018        548            999
XI93               bfr                       1017         1035         958           949         288            548
XI94               bfr                       1036         223          1035          217         224            288
XI95               bfr                       1002         274          223           1038        927            224
XI96               bfr                       1027         429          274           1019        278            927
XI97               bfr                       147          858          218           943         235            214
XI98               bfr                       247          959          858           232         230            235
XI99               bfr                       975          748          959           237         746            230
XI14               boost2_3_f3               822          728          255           529         567            538                    726   313
XI340              boost2_3_f3               790          666          728           468         539            524                    78    726
XI312              boost2_4_f4               1099         734          970           937         836            819                    797   507   272
XI313              boost2_4_f4               1100         970          1031          832         826            1000                   1047  272   1048
XI314              boost2_4_f4               771          1031         605           803         964            867                    873   1048  576
XI316              boost2_4_f4               1096         1032         206           765         744            750                    741   809   102
XI321              boost2_4_f4               1097         206          917           760         752            713                    702   102   164
XI322              boost2_4_f4               976          917          735           733         738            691                    951   164   861
XI323              boost2_4_f4               1094         370          253           1008        1012           1010                   1046  64    137
XI326              boost2_4_f4               1095         253          948           1037        1003           925                    967   137   106
XI329              boost2_4_f4               945          948          756           985         1023           898                    950   106   755
XI341              boost2_4_f4               1            731          560           944         935            916                    426   730   382
XI344              boost2_4_f4               474          560          340           386         924            909                    881   382   665
XI347              boost2_4_f4               787          340          736           895         887            405                    352   665   729
XI349              boost2_4_f4               390          812          553           342         375            781                    396   433   546
XI352              boost2_4_f4               792          553          551           446         776            465                    810   546   337
XI355              boost2_4_f4               463          551          853           330         325            319                    321   337   601
XI358              boost2_4_f4               2            942          674           301         387            407                    371   611   675
XI361              boost2_4_f4               363          674          676           394         391            451                    353   675   683
XI364              boost2_4_f4               362          676          496           356         450            308                    388   683   727
XI366              boost2_4_f4               420          687          751           310         307            393                    341   686   550
XI367              boost2_4_f4               336          597          693           417         343            466                    364   725   694
XI370              boost2_4_f4               316          693          687           379         360            438                    329   694   686
XI307              maj_bbb                   937          832          803           914         1005           976                    419   939
XI310              maj_bbb                   978          856          1020          735         11             1101                   861   602
XI315              maj_bbb                   765          760          733           663         911            945                    670   244
XI318              maj_bbb                   754          934          724           756         243            1098                   755   248
XI324              maj_bbb                   1008         1037         985           66          290            787                    67    124
XI330              maj_bbb                   989          1043         926           736         849            165                    729   289
XI342              maj_bbb                   944          386          895           15          578            463                    16    575
XI348              maj_bbb                   350          345          443           853         519            185                    601   415
XI350              maj_bbb                   342          446          330           851         685            420                    753   684
XI356              maj_bbb                   381          327          361           751         516            199                    550   606
XI357              maj_bbb                   444          434          374           496         195            205                    727   470
XI359              maj_bbb                   301          394          356           210         673            317                    1106  677
XI365              maj_bbb                   378          408          423           207         749            747                    208   202
XI372              maj_bbb                   417          379          310           464         696            362                    745   695
XI311              maj_bbi                   797          1047         873           89          298            1020                   95    1045
XI317              maj_bbi                   741          702          951           1001        960            724                    893   1025
XI328              maj_bbi                   1046         967          950           963         293            926                    991   292
XI346              maj_bbi                   426          881          352           659         428            443                    660   742
XI354              maj_bbi                   396          810          321           536         186            361                    540   430
XI363              maj_bbi                   371          353          388           682         740            423                    681   203
XI368              maj_bbi                   364          329          341           692         365            374                    690   200
XI309              maj_bib                   819          1000         867           1033        89             856                    1007  95
XI319              maj_bib                   750          713          691           280         1001           934                    276   893
XI327              maj_bib                   1010         925          898           117         963            1043                   984   991
XI345              maj_bib                   916          909          405           661         659            345                    449   660
XI353              maj_bib                   781          465          319           532         536            327                    527   540
XI362              maj_bib                   407          451          308           678         682            408                    679   681
XI369              maj_bib                   466          438          393           689         692            434                    688   690
XI308              maj_ibb                   836          826          964           1005        1033           978                    939   1007
XI320              maj_ibb                   744          752          738           911         280            754                    244   276
XI325              maj_ibb                   1012         1003         1023          290         117            989                    124   984
XI343              maj_ibb                   935          924          887           578         661            350                    575   449
XI351              maj_ibb                   375          776          325           685         532            381                    684   527
XI360              maj_ibb                   387          391          450           673         678            378                    677   679
XI371              maj_ibb                   343          360          307           696         689            444                    695   688
XI339              or_bb                     334          495          605           871         1102           576                    313
XSUM0              sink                      632          655          0             294         0
XSUM1              sink                      531          629          655           610         294
XSUM2              sink                      621          485          629           318         610
XSUM3              sink                      598          299          485           627         318
XSUM4              sink                      639          609          299           528         627
XSUM5              sink                      641          500          609           323         528
XSUM6              sink                      645          652          500           559         323
XSUM7              sink                      332          547          652           603         559
XSUM8              sink                      544          590          547           328         603
*end of top cell   8bit_RCA_ene_opt_booster


.tran              {{t_step}}ps              {{end}}ps    {{begin}}ps  {{t_step}}ps
.FiLE              {{out_file_name}}
.print             i(Rac1)
*vac1_tot
.print             nodev                     1105         0

.print             i(Rac2)
*vac2_tot
.print             nodev                     1108         0

*vac1_DUT
.print             nodev                     1104         1103
*vac2_DUT
.print             nodev                     1107         1106