.model             jjmod                jj(Rtype=1,  Vg=2.8mV,    Cap=0.064pF,  R0=100ohm,  Rn=17ohm,      Icrit=0.1mA)


.subckt            bfr                  1            2            3             12          13             14
*inst name         cell_name            a            din          dout          q           xin            xout
B1                 9                    0            jjmod        area=0.5
B2                 5                    0            jjmod        area=0.5
Kd1                Ld                   L1           -0.133
Kd2                Ld                   L2           -0.133
Kdout              Ld                   Lout         0.0
Kdq                Ld                   Lq           0.0
Kout               Lq                   Lout         -0.495
Kx1                Lx                   L1           -0.186
Kx2                Lx                   L2           -0.186
Kxd                Lx                   Ld           0.19
Kxout              Lx                   Lout         0.0
Kxq                Lx                   Lq           0.0
L1                 8                    9            1.59pH
L2                 5                    8            1.59pH
Ld                 2                    3            7.45pH
Lin                1                    8            1.23pH
Lout               6                    12           31.2pH
Lq                 8                    0            7.92pH
Lx                 13                   14           7.4pH
R1                 6                    0            1e-12ohm
.ends


.subckt            branch3              1            2            3             4
*inst name         cell_name            a            b            c             d
Lip                7                    4            0.312pH
Lp1                1                    6            11.8pH
Lp2                2                    7            10.2pH
Lp3                3                    5            11.8pH
R0                 6                    7            1e-12ohm
R1                 5                    7            1e-12ohm
.ends


.subckt            const0               1            2            11            12          13
*inst name         cell_name            din          dout         q             xin         xout
B1                 8                    0            jjmod        area=0.5
B2                 4                    0            jjmod        area=0.5
Kd1                Ld                   L1           -0.128
Kd2                Ld                   L2           -0.135
Kdout              Ld                   Lout         -0.000253
Kdq                Ld                   Lq           -0.00468
Kout               Lq                   Lout         -0.495
Kx1                Lx                   L1           -0.185
Kx2                Lx                   L2           -0.189
Kxd                Lx                   Ld           0.193
Kxout              Lx                   Lout         -7.94e-05
Kxq                Lx                   Lq           -0.00421
L1                 7                    8            1.56pH
L2                 4                    7            1.66pH
Ld                 1                    2            7.49pH
Lout               5                    11           31.2pH
Lq                 7                    0            7.82pH
Lx                 12                   13           7.47pH
R1                 5                    0            1e-12ohm
.ends


.subckt            and_bb               1            2            3             4           12             13                     14
*inst name         cell_name            a            b            din           dout        q              xin                    xout
XI0                bfr                  1            3            8             9           13             5
XI2                bfr                  2            11           4             10          7              14
XI3                branch3              9            6            10            12
XI1                const0               8            11           6             5           7
.ends


.subckt            sink                 1            2            3             10          11
*inst name         cell_name            a            din          dout          xin         xout
B1                 8                    0            jjmod        area=0.5
B2                 5                    0            jjmod        area=0.5
Kd1                Ld                   L1           -0.133
Kd2                Ld                   L2           -0.133
Kdq                Ld                   Lq           0.0
Kx1                Lx                   L1           -0.186
Kx2                Lx                   L2           -0.186
Kxd                Lx                   Ld           0.19
Kxq                Lx                   Lq           0.0
L1                 7                    8            1.59pH
L2                 5                    7            1.59pH
Ld                 2                    3            7.45pH
Lin                1                    7            1.23pH
Lq                 7                    0            7.92pH
Lx                 10                   11           7.4pH
.ends


*this is top cell  and2_hstp033_energy
R1                 9                    48           1000.0ohm
R3                 10                   46           1000.0ohm
R9                 6                    34           100000.0ohm
Rac1               7                    52           100000.0ohm
Rac2               4                    19           100000.0ohm
V1                 9                    0            PWL          (0ps          0mv         20ps           {{input[0]}})
V3                 10                   0            PWL          (0ps          0mv         20ps           {{input[1]}})
VDC                6                    0            PWL          (0ps          0mV         20ps           113000mV)
V0                 7                    0            SIN          (0            81000mV     {{freq}}MEGHz  {{40+period|int/4}}ps  0)
V2                 4                    0            SIN          (0            81000mV     {{freq}}MEGHz  40ps                   0)
XI20               and_bb               17           13           47            49          29             51                     50
XI1                bfr                  48           34           31            28          52             33
XI10               bfr                  27           18           36            45          51             35
XI12               bfr                  21           36           12            14          35             26
XI14               bfr                  45           47           38            17          32             11
XI16               bfr                  14           38           12            13          11             20
XI21               bfr                  30           39           44            24          43             50
XI23               bfr                  24           42           44            23          0              37
XI24               bfr                  29           39           49            30          32             37
XI3                bfr                  46           31           25            22          33             26
XI5                bfr                  28           18           16            27          19             15
XI7                bfr                  22           16           25            21          15             20
XI22               sink                 23           42           0             43          0
*end of top cell   and2_hstp033_energy


.tran              {{t_step}}ps         {{end}}ps    {{begin}}ps  {{t_step}}ps
.FiLE              {{out_file_name}}
.print             i(Rac1)
*vac1_tot
.print             nodev                52           0

.print             i(Rac2)
*vac1_DUT
.print             nodev                51           50